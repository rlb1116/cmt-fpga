-- fpacc64.vhd

-- Generated using ACDS version 16.0 211

library IEEE;
library altera_fp_acc_custom_160;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity fpacc64 is
	port (
		ao     : out std_logic;                                        --     ao.ao
		areset : in  std_logic                     := '0';             -- areset.reset
		clk    : in  std_logic                     := '0';             --    clk.clk
		en     : in  std_logic_vector(0 downto 0)  := (others => '0'); --     en.en
		n      : in  std_logic                     := '0';             --      n.n
		r      : out std_logic_vector(63 downto 0);                    --      r.r
		x      : in  std_logic_vector(63 downto 0) := (others => '0'); --      x.x
		xo     : out std_logic;                                        --     xo.xo
		xu     : out std_logic                                         --     xu.xu
	);
end entity fpacc64;

architecture rtl of fpacc64 is
	component fpacc64_altera_fp_acc_custom_160_bhzzlly is
		port (
			clk    : in  std_logic                     := 'X';             -- clk
			areset : in  std_logic                     := 'X';             -- reset
			x      : in  std_logic_vector(63 downto 0) := (others => 'X'); -- x
			n      : in  std_logic                     := 'X';             -- n
			r      : out std_logic_vector(63 downto 0);                    -- r
			xo     : out std_logic;                                        -- xo
			xu     : out std_logic;                                        -- xu
			ao     : out std_logic;                                        -- ao
			en     : in  std_logic_vector(0 downto 0)  := (others => 'X')  -- en
		);
	end component fpacc64_altera_fp_acc_custom_160_bhzzlly;

	for fp_acc_custom_0 : fpacc64_altera_fp_acc_custom_160_bhzzlly
		use entity altera_fp_acc_custom_160.fpacc64_altera_fp_acc_custom_160_bhzzlly;
begin

	fp_acc_custom_0 : component fpacc64_altera_fp_acc_custom_160_bhzzlly
		port map (
			clk    => clk,    --    clk.clk
			areset => areset, -- areset.reset
			x      => x,      --      x.x
			n      => n,      --      n.n
			r      => r,      --      r.r
			xo     => xo,     --     xo.xo
			xu     => xu,     --     xu.xu
			ao     => ao,     --     ao.ao
			en     => en      --     en.en
		);

end architecture rtl; -- of fpacc64
