// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, the Altera Quartus Prime License Agreement,
// the Altera MegaCore Function License Agreement, or other 
// applicable license agreement, including, without limitation, 
// that your use is for the sole purpose of programming logic 
// devices manufactured by Altera and sold by Altera or its 
// authorized distributors.  Please refer to the applicable 
// agreement for further details.

// VENDOR "Altera"
// PROGRAM "Quartus Prime"
// VERSION "Version 16.0.0 Build 211 04/27/2016 SJ Pro Edition"

// DATE "03/26/2019 17:07:55"

// 
// Device: Altera 10AX048E1F29E1SG Package FBGA780
// 

// 
// This greybox netlist file is for third party Synthesis Tools
// for timing and resource estimation only.
// 


module fpmult64 (
	q,
	clk,
	areset,
	en,
	b,
	a)/* synthesis synthesis_greybox=0 */;
output 	[63:0] q;
input 	clk;
input 	areset;
input 	[0:0] en;
input 	[63:0] b;
input 	[63:0] a;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \fp_functions_0|add_7~1_sumout ;
wire \fp_functions_0|add_8~1_sumout ;
wire \fp_functions_0|add_6~1_sumout ;
wire \fp_functions_0|add_6~2 ;
wire \fp_functions_0|add_7~6_cout ;
wire \fp_functions_0|add_8~6_cout ;
wire \fp_functions_0|add_6~5_sumout ;
wire \fp_functions_0|add_6~6 ;
wire \fp_functions_0|add_6~9_sumout ;
wire \fp_functions_0|add_6~10 ;
wire \fp_functions_0|add_6~13_sumout ;
wire \fp_functions_0|add_6~14 ;
wire \fp_functions_0|add_6~17_sumout ;
wire \fp_functions_0|add_6~18 ;
wire \fp_functions_0|add_6~21_sumout ;
wire \fp_functions_0|add_6~22 ;
wire \fp_functions_0|add_6~25_sumout ;
wire \fp_functions_0|add_6~26 ;
wire \fp_functions_0|add_6~29_sumout ;
wire \fp_functions_0|add_6~30 ;
wire \fp_functions_0|add_6~33_sumout ;
wire \fp_functions_0|add_6~34 ;
wire \fp_functions_0|add_6~37_sumout ;
wire \fp_functions_0|add_6~38 ;
wire \fp_functions_0|add_6~41_sumout ;
wire \fp_functions_0|add_6~42 ;
wire \fp_functions_0|add_6~45_sumout ;
wire \fp_functions_0|add_6~46 ;
wire \fp_functions_0|add_6~49_sumout ;
wire \fp_functions_0|add_6~50 ;
wire \fp_functions_0|add_6~53_sumout ;
wire \fp_functions_0|add_6~54 ;
wire \fp_functions_0|add_6~57_sumout ;
wire \fp_functions_0|add_6~58 ;
wire \fp_functions_0|add_6~61_sumout ;
wire \fp_functions_0|add_6~62 ;
wire \fp_functions_0|add_6~65_sumout ;
wire \fp_functions_0|add_6~66 ;
wire \fp_functions_0|add_6~69_sumout ;
wire \fp_functions_0|add_6~70 ;
wire \fp_functions_0|add_6~73_sumout ;
wire \fp_functions_0|add_6~74 ;
wire \fp_functions_0|add_6~77_sumout ;
wire \fp_functions_0|add_6~78 ;
wire \fp_functions_0|add_6~81_sumout ;
wire \fp_functions_0|add_6~82 ;
wire \fp_functions_0|add_6~85_sumout ;
wire \fp_functions_0|add_6~86 ;
wire \fp_functions_0|add_6~89_sumout ;
wire \fp_functions_0|add_6~90 ;
wire \fp_functions_0|add_6~93_sumout ;
wire \fp_functions_0|add_6~94 ;
wire \fp_functions_0|add_6~97_sumout ;
wire \fp_functions_0|add_6~98 ;
wire \fp_functions_0|add_6~101_sumout ;
wire \fp_functions_0|add_6~102 ;
wire \fp_functions_0|add_6~105_sumout ;
wire \fp_functions_0|add_6~106 ;
wire \fp_functions_0|add_6~109_sumout ;
wire \fp_functions_0|add_6~110 ;
wire \fp_functions_0|add_6~113_sumout ;
wire \fp_functions_0|add_6~114 ;
wire \fp_functions_0|add_6~117_sumout ;
wire \fp_functions_0|add_6~118 ;
wire \fp_functions_0|add_6~121_sumout ;
wire \fp_functions_0|add_6~122 ;
wire \fp_functions_0|add_6~125_sumout ;
wire \fp_functions_0|add_6~126 ;
wire \fp_functions_0|add_6~129_sumout ;
wire \fp_functions_0|add_6~130 ;
wire \fp_functions_0|add_6~133_sumout ;
wire \fp_functions_0|add_6~134 ;
wire \fp_functions_0|add_6~137_sumout ;
wire \fp_functions_0|add_6~138 ;
wire \fp_functions_0|add_6~141_sumout ;
wire \fp_functions_0|add_6~142 ;
wire \fp_functions_0|add_6~145_sumout ;
wire \fp_functions_0|add_6~146 ;
wire \fp_functions_0|add_6~149_sumout ;
wire \fp_functions_0|add_6~150 ;
wire \fp_functions_0|add_6~153_sumout ;
wire \fp_functions_0|add_6~154 ;
wire \fp_functions_0|add_6~157_sumout ;
wire \fp_functions_0|add_6~158 ;
wire \fp_functions_0|add_6~161_sumout ;
wire \fp_functions_0|add_6~162 ;
wire \fp_functions_0|add_6~165_sumout ;
wire \fp_functions_0|add_6~166 ;
wire \fp_functions_0|add_6~169_sumout ;
wire \fp_functions_0|add_6~170 ;
wire \fp_functions_0|add_6~173_sumout ;
wire \fp_functions_0|add_6~174 ;
wire \fp_functions_0|add_6~177_sumout ;
wire \fp_functions_0|add_6~178 ;
wire \fp_functions_0|add_6~181_sumout ;
wire \fp_functions_0|add_6~182 ;
wire \fp_functions_0|add_6~185_sumout ;
wire \fp_functions_0|add_6~186 ;
wire \fp_functions_0|add_6~189_sumout ;
wire \fp_functions_0|add_6~190 ;
wire \fp_functions_0|add_6~193_sumout ;
wire \fp_functions_0|add_6~194 ;
wire \fp_functions_0|add_6~197_sumout ;
wire \fp_functions_0|add_6~198 ;
wire \fp_functions_0|add_6~201_sumout ;
wire \fp_functions_0|add_6~202 ;
wire \fp_functions_0|add_6~205_sumout ;
wire \fp_functions_0|add_6~206 ;
wire \fp_functions_0|add_6~209_sumout ;
wire \fp_functions_0|add_6~210 ;
wire \fp_functions_0|add_6~213_sumout ;
wire \fp_functions_0|add_6~214 ;
wire \fp_functions_0|add_6~217_sumout ;
wire \fp_functions_0|add_6~218 ;
wire \fp_functions_0|add_6~221_sumout ;
wire \fp_functions_0|add_6~222 ;
wire \fp_functions_0|add_6~225_sumout ;
wire \fp_functions_0|add_6~226 ;
wire \fp_functions_0|add_6~229_sumout ;
wire \fp_functions_0|add_6~230 ;
wire \fp_functions_0|add_6~233_sumout ;
wire \fp_functions_0|add_6~234 ;
wire \fp_functions_0|add_6~237_sumout ;
wire \fp_functions_0|add_6~238 ;
wire \fp_functions_0|add_6~241_sumout ;
wire \fp_functions_0|add_6~242 ;
wire \fp_functions_0|add_6~245_sumout ;
wire \fp_functions_0|add_6~246 ;
wire \fp_functions_0|add_6~249_sumout ;
wire \fp_functions_0|add_6~250 ;
wire \fp_functions_0|add_6~254_cout ;
wire \fp_functions_0|add_6~257_sumout ;
wire \fp_functions_0|add_7~10_cout ;
wire \fp_functions_0|add_8~10_cout ;
wire \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[1]~q ;
wire \fp_functions_0|add_6~261_sumout ;
wire \fp_functions_0|add_6~262 ;
wire \fp_functions_0|add_7~14_cout ;
wire \fp_functions_0|add_8~14_cout ;
wire \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[2]~q ;
wire \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[3]~q ;
wire \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[4]~q ;
wire \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[5]~q ;
wire \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[6]~q ;
wire \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[7]~q ;
wire \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[8]~q ;
wire \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[9]~q ;
wire \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[10]~q ;
wire \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[11]~q ;
wire \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[12]~q ;
wire \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[13]~q ;
wire \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[14]~q ;
wire \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[15]~q ;
wire \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[16]~q ;
wire \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[17]~q ;
wire \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[18]~q ;
wire \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[19]~q ;
wire \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[20]~q ;
wire \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[21]~q ;
wire \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[22]~q ;
wire \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[23]~q ;
wire \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[24]~q ;
wire \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[25]~q ;
wire \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[26]~q ;
wire \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[27]~q ;
wire \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[28]~q ;
wire \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[29]~q ;
wire \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[30]~q ;
wire \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[31]~q ;
wire \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[32]~q ;
wire \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[33]~q ;
wire \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[34]~q ;
wire \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[35]~q ;
wire \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[36]~q ;
wire \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[37]~q ;
wire \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[38]~q ;
wire \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[39]~q ;
wire \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[40]~q ;
wire \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[41]~q ;
wire \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[42]~q ;
wire \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[43]~q ;
wire \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[44]~q ;
wire \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[45]~q ;
wire \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[46]~q ;
wire \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[47]~q ;
wire \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[48]~q ;
wire \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[49]~q ;
wire \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[50]~q ;
wire \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[51]~q ;
wire \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[52]~q ;
wire \fp_functions_0|add_5~1_sumout ;
wire \fp_functions_0|add_5~2 ;
wire \fp_functions_0|add_5~5_sumout ;
wire \fp_functions_0|add_5~6 ;
wire \fp_functions_0|add_5~9_sumout ;
wire \fp_functions_0|add_5~10 ;
wire \fp_functions_0|add_5~13_sumout ;
wire \fp_functions_0|add_5~14 ;
wire \fp_functions_0|add_5~17_sumout ;
wire \fp_functions_0|add_5~18 ;
wire \fp_functions_0|add_5~21_sumout ;
wire \fp_functions_0|add_5~22 ;
wire \fp_functions_0|add_5~25_sumout ;
wire \fp_functions_0|add_5~26 ;
wire \fp_functions_0|add_5~29_sumout ;
wire \fp_functions_0|add_5~30 ;
wire \fp_functions_0|add_5~33_sumout ;
wire \fp_functions_0|add_5~34 ;
wire \fp_functions_0|add_5~37_sumout ;
wire \fp_functions_0|add_5~38 ;
wire \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[0]~q ;
wire \fp_functions_0|add_5~41_sumout ;
wire \fp_functions_0|add_6~265_sumout ;
wire \fp_functions_0|add_6~266 ;
wire \fp_functions_0|add_7~18_cout ;
wire \fp_functions_0|add_8~18_cout ;
wire \fp_functions_0|add_1~1_sumout ;
wire \fp_functions_0|add_1~2 ;
wire \fp_functions_0|add_1~5_sumout ;
wire \fp_functions_0|add_1~6 ;
wire \fp_functions_0|add_1~9_sumout ;
wire \fp_functions_0|add_5~45_sumout ;
wire \fp_functions_0|add_5~46 ;
wire \fp_functions_0|add_6~269_sumout ;
wire \fp_functions_0|add_6~270 ;
wire \fp_functions_0|add_7~22_cout ;
wire \fp_functions_0|add_8~22_cout ;
wire \fp_functions_0|add_1~13_sumout ;
wire \fp_functions_0|add_1~14 ;
wire \fp_functions_0|add_1~17_sumout ;
wire \fp_functions_0|add_1~18 ;
wire \fp_functions_0|add_1~21_sumout ;
wire \fp_functions_0|add_1~22 ;
wire \fp_functions_0|add_1~25_sumout ;
wire \fp_functions_0|add_1~26 ;
wire \fp_functions_0|add_1~29_sumout ;
wire \fp_functions_0|add_1~30 ;
wire \fp_functions_0|add_1~33_sumout ;
wire \fp_functions_0|add_1~34 ;
wire \fp_functions_0|add_1~37_sumout ;
wire \fp_functions_0|add_1~38 ;
wire \fp_functions_0|add_1~41_sumout ;
wire \fp_functions_0|add_1~42 ;
wire \fp_functions_0|add_1~45_sumout ;
wire \fp_functions_0|add_1~46 ;
wire \fp_functions_0|add_1~49_sumout ;
wire \fp_functions_0|add_1~50 ;
wire \fp_functions_0|add_1~53_sumout ;
wire \fp_functions_0|add_1~54 ;
wire \fp_functions_0|add_1~57_sumout ;
wire \fp_functions_0|add_1~58 ;
wire \fp_functions_0|add_1~61_sumout ;
wire \fp_functions_0|add_1~62 ;
wire \fp_functions_0|add_1~65_sumout ;
wire \fp_functions_0|add_1~66 ;
wire \fp_functions_0|add_1~69_sumout ;
wire \fp_functions_0|add_1~70 ;
wire \fp_functions_0|add_1~73_sumout ;
wire \fp_functions_0|add_1~74 ;
wire \fp_functions_0|add_1~77_sumout ;
wire \fp_functions_0|add_1~78 ;
wire \fp_functions_0|add_1~81_sumout ;
wire \fp_functions_0|add_1~82 ;
wire \fp_functions_0|add_1~85_sumout ;
wire \fp_functions_0|add_1~86 ;
wire \fp_functions_0|add_1~89_sumout ;
wire \fp_functions_0|add_1~90 ;
wire \fp_functions_0|add_1~93_sumout ;
wire \fp_functions_0|add_1~94 ;
wire \fp_functions_0|add_1~97_sumout ;
wire \fp_functions_0|add_1~98 ;
wire \fp_functions_0|add_1~101_sumout ;
wire \fp_functions_0|add_1~102 ;
wire \fp_functions_0|add_1~105_sumout ;
wire \fp_functions_0|add_1~106 ;
wire \fp_functions_0|add_1~109_sumout ;
wire \fp_functions_0|add_1~110 ;
wire \fp_functions_0|add_1~113_sumout ;
wire \fp_functions_0|add_1~114 ;
wire \fp_functions_0|add_1~117_sumout ;
wire \fp_functions_0|add_1~118 ;
wire \fp_functions_0|add_1~121_sumout ;
wire \fp_functions_0|add_1~122 ;
wire \fp_functions_0|add_1~125_sumout ;
wire \fp_functions_0|add_1~126 ;
wire \fp_functions_0|add_1~129_sumout ;
wire \fp_functions_0|add_1~130 ;
wire \fp_functions_0|add_1~133_sumout ;
wire \fp_functions_0|add_1~134 ;
wire \fp_functions_0|add_1~137_sumout ;
wire \fp_functions_0|add_1~138 ;
wire \fp_functions_0|add_1~141_sumout ;
wire \fp_functions_0|add_1~142 ;
wire \fp_functions_0|add_1~145_sumout ;
wire \fp_functions_0|add_1~146 ;
wire \fp_functions_0|add_1~149_sumout ;
wire \fp_functions_0|add_1~150 ;
wire \fp_functions_0|add_1~153_sumout ;
wire \fp_functions_0|add_1~154 ;
wire \fp_functions_0|add_1~157_sumout ;
wire \fp_functions_0|add_1~158 ;
wire \fp_functions_0|add_1~161_sumout ;
wire \fp_functions_0|add_1~162 ;
wire \fp_functions_0|add_1~165_sumout ;
wire \fp_functions_0|add_1~166 ;
wire \fp_functions_0|add_1~169_sumout ;
wire \fp_functions_0|add_1~170 ;
wire \fp_functions_0|add_1~173_sumout ;
wire \fp_functions_0|add_1~174 ;
wire \fp_functions_0|add_1~177_sumout ;
wire \fp_functions_0|add_1~178 ;
wire \fp_functions_0|add_1~181_sumout ;
wire \fp_functions_0|add_1~182 ;
wire \fp_functions_0|add_1~185_sumout ;
wire \fp_functions_0|add_1~186 ;
wire \fp_functions_0|add_1~189_sumout ;
wire \fp_functions_0|add_1~190 ;
wire \fp_functions_0|add_1~193_sumout ;
wire \fp_functions_0|add_1~194 ;
wire \fp_functions_0|add_1~197_sumout ;
wire \fp_functions_0|add_1~198 ;
wire \fp_functions_0|add_1~201_sumout ;
wire \fp_functions_0|add_1~202 ;
wire \fp_functions_0|add_1~205_sumout ;
wire \fp_functions_0|add_1~206 ;
wire \fp_functions_0|add_1~209_sumout ;
wire \fp_functions_0|add_1~210 ;
wire \fp_functions_0|add_1~213_sumout ;
wire \fp_functions_0|add_1~214 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_wire[0] ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0~PORTBDATAOUT1 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0~PORTBDATAOUT2 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0~PORTBDATAOUT3 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0~PORTBDATAOUT4 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0~PORTBDATAOUT5 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0~PORTBDATAOUT6 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0~PORTBDATAOUT7 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0~PORTBDATAOUT8 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0~PORTBDATAOUT9 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0~PORTBDATAOUT10 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0~PORTBDATAOUT11 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0~PORTBDATAOUT12 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0~PORTBDATAOUT13 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0~PORTBDATAOUT14 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0~PORTBDATAOUT15 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0~PORTBDATAOUT16 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0~PORTBDATAOUT17 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0~PORTBDATAOUT18 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0~PORTBDATAOUT19 ;
wire \fp_functions_0|add_1~217_sumout ;
wire \fp_functions_0|add_1~218 ;
wire \fp_functions_0|add_1~221_sumout ;
wire \fp_functions_0|add_1~222 ;
wire \fp_functions_0|add_1~225_sumout ;
wire \fp_functions_0|add_1~226 ;
wire \fp_functions_0|add_1~229_sumout ;
wire \fp_functions_0|add_1~230 ;
wire \fp_functions_0|add_1~233_sumout ;
wire \fp_functions_0|add_1~234 ;
wire \fp_functions_0|add_1~237_sumout ;
wire \fp_functions_0|add_1~238 ;
wire \fp_functions_0|add_1~241_sumout ;
wire \fp_functions_0|add_1~242 ;
wire \fp_functions_0|add_1~245_sumout ;
wire \fp_functions_0|add_1~246 ;
wire \fp_functions_0|add_1~249_sumout ;
wire \fp_functions_0|add_1~250 ;
wire \fp_functions_0|add_1~253_sumout ;
wire \fp_functions_0|add_1~254 ;
wire \fp_functions_0|add_1~257_sumout ;
wire \fp_functions_0|add_1~258 ;
wire \fp_functions_0|add_1~261_sumout ;
wire \fp_functions_0|add_1~262 ;
wire \fp_functions_0|add_1~265_sumout ;
wire \fp_functions_0|add_1~266 ;
wire \fp_functions_0|add_1~269_sumout ;
wire \fp_functions_0|add_1~270 ;
wire \fp_functions_0|add_1~273_sumout ;
wire \fp_functions_0|add_1~274 ;
wire \fp_functions_0|add_1~277_sumout ;
wire \fp_functions_0|add_1~278 ;
wire \fp_functions_0|add_1~281_sumout ;
wire \fp_functions_0|add_1~282 ;
wire \fp_functions_0|add_1~285_sumout ;
wire \fp_functions_0|add_1~286 ;
wire \fp_functions_0|add_1~289_sumout ;
wire \fp_functions_0|add_1~290 ;
wire \fp_functions_0|add_1~293_sumout ;
wire \fp_functions_0|add_1~294 ;
wire \fp_functions_0|add_1~297_sumout ;
wire \fp_functions_0|add_1~298 ;
wire \fp_functions_0|add_1~301_sumout ;
wire \fp_functions_0|add_1~302 ;
wire \fp_functions_0|add_1~305_sumout ;
wire \fp_functions_0|add_1~306 ;
wire \fp_functions_0|add_1~309_sumout ;
wire \fp_functions_0|add_1~310 ;
wire \fp_functions_0|add_1~313_sumout ;
wire \fp_functions_0|add_1~314 ;
wire \fp_functions_0|add_1~317_sumout ;
wire \fp_functions_0|add_1~318 ;
wire \fp_functions_0|add_1~321_sumout ;
wire \fp_functions_0|add_1~322 ;
wire \fp_functions_0|add_5~49_sumout ;
wire \fp_functions_0|add_5~50 ;
wire \fp_functions_0|add_7~26_cout ;
wire \fp_functions_0|add_8~26_cout ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_wire[1] ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1~PORTBDATAOUT1 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1~PORTBDATAOUT2 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1~PORTBDATAOUT3 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1~PORTBDATAOUT4 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1~PORTBDATAOUT5 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1~PORTBDATAOUT6 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1~PORTBDATAOUT7 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1~PORTBDATAOUT8 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1~PORTBDATAOUT9 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1~PORTBDATAOUT10 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1~PORTBDATAOUT11 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1~PORTBDATAOUT12 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1~PORTBDATAOUT13 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1~PORTBDATAOUT14 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1~PORTBDATAOUT15 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1~PORTBDATAOUT16 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1~PORTBDATAOUT17 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1~PORTBDATAOUT18 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1~PORTBDATAOUT19 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_wire[2] ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2~PORTBDATAOUT1 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2~PORTBDATAOUT2 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2~PORTBDATAOUT3 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2~PORTBDATAOUT4 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2~PORTBDATAOUT5 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2~PORTBDATAOUT6 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2~PORTBDATAOUT7 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2~PORTBDATAOUT8 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2~PORTBDATAOUT9 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2~PORTBDATAOUT10 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2~PORTBDATAOUT11 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2~PORTBDATAOUT12 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2~PORTBDATAOUT13 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2~PORTBDATAOUT14 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2~PORTBDATAOUT15 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2~PORTBDATAOUT16 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2~PORTBDATAOUT17 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2~PORTBDATAOUT18 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2~PORTBDATAOUT19 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_wire[3] ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3~PORTBDATAOUT1 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3~PORTBDATAOUT2 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3~PORTBDATAOUT3 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3~PORTBDATAOUT4 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3~PORTBDATAOUT5 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3~PORTBDATAOUT6 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3~PORTBDATAOUT7 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3~PORTBDATAOUT8 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3~PORTBDATAOUT9 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3~PORTBDATAOUT10 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3~PORTBDATAOUT11 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3~PORTBDATAOUT12 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3~PORTBDATAOUT13 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3~PORTBDATAOUT14 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3~PORTBDATAOUT15 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3~PORTBDATAOUT16 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3~PORTBDATAOUT17 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3~PORTBDATAOUT18 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3~PORTBDATAOUT19 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_wire[4] ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4~PORTBDATAOUT1 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4~PORTBDATAOUT2 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4~PORTBDATAOUT3 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4~PORTBDATAOUT4 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4~PORTBDATAOUT5 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4~PORTBDATAOUT6 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4~PORTBDATAOUT7 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4~PORTBDATAOUT8 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4~PORTBDATAOUT9 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4~PORTBDATAOUT10 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4~PORTBDATAOUT11 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4~PORTBDATAOUT12 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4~PORTBDATAOUT13 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4~PORTBDATAOUT14 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4~PORTBDATAOUT15 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4~PORTBDATAOUT16 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4~PORTBDATAOUT17 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4~PORTBDATAOUT18 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4~PORTBDATAOUT19 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_wire[5] ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5~PORTBDATAOUT1 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5~PORTBDATAOUT2 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5~PORTBDATAOUT3 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5~PORTBDATAOUT4 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5~PORTBDATAOUT5 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5~PORTBDATAOUT6 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5~PORTBDATAOUT7 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5~PORTBDATAOUT8 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5~PORTBDATAOUT9 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5~PORTBDATAOUT10 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5~PORTBDATAOUT11 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5~PORTBDATAOUT12 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5~PORTBDATAOUT13 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5~PORTBDATAOUT14 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5~PORTBDATAOUT15 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5~PORTBDATAOUT16 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5~PORTBDATAOUT17 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5~PORTBDATAOUT18 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5~PORTBDATAOUT19 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_wire[6] ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6~PORTBDATAOUT1 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6~PORTBDATAOUT2 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6~PORTBDATAOUT3 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6~PORTBDATAOUT4 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6~PORTBDATAOUT5 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6~PORTBDATAOUT6 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6~PORTBDATAOUT7 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6~PORTBDATAOUT8 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6~PORTBDATAOUT9 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6~PORTBDATAOUT10 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6~PORTBDATAOUT11 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6~PORTBDATAOUT12 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6~PORTBDATAOUT13 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6~PORTBDATAOUT14 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6~PORTBDATAOUT15 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6~PORTBDATAOUT16 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6~PORTBDATAOUT17 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6~PORTBDATAOUT18 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6~PORTBDATAOUT19 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_wire[7] ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7~PORTBDATAOUT1 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7~PORTBDATAOUT2 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7~PORTBDATAOUT3 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7~PORTBDATAOUT4 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7~PORTBDATAOUT5 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7~PORTBDATAOUT6 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7~PORTBDATAOUT7 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7~PORTBDATAOUT8 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7~PORTBDATAOUT9 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7~PORTBDATAOUT10 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7~PORTBDATAOUT11 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7~PORTBDATAOUT12 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7~PORTBDATAOUT13 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7~PORTBDATAOUT14 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7~PORTBDATAOUT15 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7~PORTBDATAOUT16 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7~PORTBDATAOUT17 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7~PORTBDATAOUT18 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7~PORTBDATAOUT19 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_wire[8] ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8~PORTBDATAOUT1 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8~PORTBDATAOUT2 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8~PORTBDATAOUT3 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8~PORTBDATAOUT4 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8~PORTBDATAOUT5 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8~PORTBDATAOUT6 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8~PORTBDATAOUT7 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8~PORTBDATAOUT8 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8~PORTBDATAOUT9 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8~PORTBDATAOUT10 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8~PORTBDATAOUT11 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8~PORTBDATAOUT12 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8~PORTBDATAOUT13 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8~PORTBDATAOUT14 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8~PORTBDATAOUT15 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8~PORTBDATAOUT16 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8~PORTBDATAOUT17 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8~PORTBDATAOUT18 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8~PORTBDATAOUT19 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_wire[9] ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9~PORTBDATAOUT1 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9~PORTBDATAOUT2 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9~PORTBDATAOUT3 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9~PORTBDATAOUT4 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9~PORTBDATAOUT5 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9~PORTBDATAOUT6 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9~PORTBDATAOUT7 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9~PORTBDATAOUT8 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9~PORTBDATAOUT9 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9~PORTBDATAOUT10 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9~PORTBDATAOUT11 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9~PORTBDATAOUT12 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9~PORTBDATAOUT13 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9~PORTBDATAOUT14 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9~PORTBDATAOUT15 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9~PORTBDATAOUT16 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9~PORTBDATAOUT17 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9~PORTBDATAOUT18 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9~PORTBDATAOUT19 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_wire[10] ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10~PORTBDATAOUT1 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10~PORTBDATAOUT2 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10~PORTBDATAOUT3 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10~PORTBDATAOUT4 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10~PORTBDATAOUT5 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10~PORTBDATAOUT6 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10~PORTBDATAOUT7 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10~PORTBDATAOUT8 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10~PORTBDATAOUT9 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10~PORTBDATAOUT10 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10~PORTBDATAOUT11 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10~PORTBDATAOUT12 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10~PORTBDATAOUT13 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10~PORTBDATAOUT14 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10~PORTBDATAOUT15 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10~PORTBDATAOUT16 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10~PORTBDATAOUT17 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10~PORTBDATAOUT18 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10~PORTBDATAOUT19 ;
wire \fp_functions_0|add_7~30_cout ;
wire \fp_functions_0|add_8~30_cout ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][0] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][1] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][2] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][3] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][4] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][5] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][6] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][7] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][8] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][9] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][10] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][11] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][12] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][13] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][14] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][15] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][16] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][17] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][18] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][19] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][20] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][21] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][22] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][23] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][24] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][25] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][26] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][27] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][28] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][29] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][30] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][31] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][32] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][33] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][34] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][35] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][36] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][37] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][38] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][39] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][40] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][41] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][42] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][43] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][44] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][45] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][46] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][47] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][48] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][49] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][50] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][51] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][52] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][53] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][54] ;
wire \fp_functions_0|mult_2~12 ;
wire \fp_functions_0|mult_2~13 ;
wire \fp_functions_0|mult_2~14 ;
wire \fp_functions_0|mult_2~15 ;
wire \fp_functions_0|mult_2~16 ;
wire \fp_functions_0|mult_2~17 ;
wire \fp_functions_0|mult_2~18 ;
wire \fp_functions_0|mult_2~19 ;
wire \fp_functions_0|mult_2~20 ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][0] ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][1] ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][2] ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][3] ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][4] ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][5] ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][6] ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][7] ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][8] ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][9] ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][10] ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][11] ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][12] ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][13] ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][14] ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][15] ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][16] ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][17] ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][18] ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][19] ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][20] ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][21] ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][22] ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][23] ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][24] ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][25] ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][26] ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][27] ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][28] ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][29] ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][30] ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][31] ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][32] ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][33] ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][34] ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][35] ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][36] ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][37] ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][38] ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][39] ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][40] ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][41] ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][42] ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][43] ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][44] ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][45] ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][46] ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][47] ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][48] ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][49] ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][50] ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][51] ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][52] ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][53] ;
wire \fp_functions_0|mult_0~12 ;
wire \fp_functions_0|mult_0~13 ;
wire \fp_functions_0|mult_0~14 ;
wire \fp_functions_0|mult_0~15 ;
wire \fp_functions_0|mult_0~16 ;
wire \fp_functions_0|mult_0~17 ;
wire \fp_functions_0|mult_0~18 ;
wire \fp_functions_0|mult_0~19 ;
wire \fp_functions_0|mult_0~20 ;
wire \fp_functions_0|mult_0~21 ;
wire \fp_functions_0|mult_1~12_resulta ;
wire \fp_functions_0|mult_1~13 ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][2] ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][3] ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][4] ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][5] ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][6] ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][7] ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][8] ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][9] ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][10] ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][11] ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][12] ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][13] ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][14] ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][15] ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][16] ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][17] ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][18] ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][19] ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][20] ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][21] ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][22] ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][23] ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][24] ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][25] ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][26] ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][27] ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][28] ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][29] ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][30] ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][31] ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][32] ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][33] ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][34] ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][35] ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][36] ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][37] ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][38] ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][39] ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][40] ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][41] ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][42] ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][43] ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][44] ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][45] ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][46] ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][47] ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][48] ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][49] ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][50] ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][51] ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][52] ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][53] ;
wire \fp_functions_0|mult_1~14 ;
wire \fp_functions_0|mult_1~15 ;
wire \fp_functions_0|mult_1~16 ;
wire \fp_functions_0|mult_1~17 ;
wire \fp_functions_0|mult_1~18 ;
wire \fp_functions_0|mult_1~19 ;
wire \fp_functions_0|mult_1~20 ;
wire \fp_functions_0|mult_1~21 ;
wire \fp_functions_0|mult_1~22 ;
wire \fp_functions_0|mult_1~23 ;
wire \fp_functions_0|add_7~34_cout ;
wire \fp_functions_0|add_8~34_cout ;
wire \fp_functions_0|add_4~1_sumout ;
wire \fp_functions_0|add_4~2 ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][0] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][1] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][2] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][3] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][4] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][5] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][6] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][7] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][8] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][9] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][10] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][11] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][12] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][13] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][14] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][15] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][16] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][17] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][18] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][19] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][20] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][21] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][22] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][23] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][24] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][25] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][26] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][27] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][28] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][29] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][30] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][31] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][32] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][33] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][34] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][35] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][36] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][37] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][38] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][39] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][40] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][41] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][42] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][43] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][44] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][45] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][46] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][47] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][48] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][49] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][50] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][51] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][52] ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][53] ;
wire \fp_functions_0|mult_3~12 ;
wire \fp_functions_0|mult_3~13 ;
wire \fp_functions_0|mult_3~14 ;
wire \fp_functions_0|mult_3~15 ;
wire \fp_functions_0|mult_3~16 ;
wire \fp_functions_0|mult_3~17 ;
wire \fp_functions_0|mult_3~18 ;
wire \fp_functions_0|mult_3~19 ;
wire \fp_functions_0|mult_3~20 ;
wire \fp_functions_0|mult_3~21 ;
wire \fp_functions_0|mult_3~86 ;
wire \fp_functions_0|mult_3~87 ;
wire \fp_functions_0|mult_3~88 ;
wire \fp_functions_0|mult_3~89 ;
wire \fp_functions_0|mult_3~90 ;
wire \fp_functions_0|mult_3~91 ;
wire \fp_functions_0|mult_3~92 ;
wire \fp_functions_0|mult_3~93 ;
wire \fp_functions_0|mult_3~94 ;
wire \fp_functions_0|mult_3~95 ;
wire \fp_functions_0|mult_3~96 ;
wire \fp_functions_0|mult_3~97 ;
wire \fp_functions_0|mult_3~98 ;
wire \fp_functions_0|mult_3~99 ;
wire \fp_functions_0|mult_3~100 ;
wire \fp_functions_0|mult_3~101 ;
wire \fp_functions_0|mult_3~102 ;
wire \fp_functions_0|mult_3~103 ;
wire \fp_functions_0|mult_3~104 ;
wire \fp_functions_0|mult_3~105 ;
wire \fp_functions_0|mult_3~106 ;
wire \fp_functions_0|mult_3~107 ;
wire \fp_functions_0|mult_3~108 ;
wire \fp_functions_0|mult_3~109 ;
wire \fp_functions_0|mult_3~110 ;
wire \fp_functions_0|mult_3~111 ;
wire \fp_functions_0|mult_3~112 ;
wire \fp_functions_0|mult_3~113 ;
wire \fp_functions_0|mult_3~114 ;
wire \fp_functions_0|mult_3~115 ;
wire \fp_functions_0|mult_3~116 ;
wire \fp_functions_0|mult_3~117 ;
wire \fp_functions_0|mult_3~118 ;
wire \fp_functions_0|mult_3~119 ;
wire \fp_functions_0|mult_3~120 ;
wire \fp_functions_0|mult_3~121 ;
wire \fp_functions_0|mult_3~122 ;
wire \fp_functions_0|mult_3~123 ;
wire \fp_functions_0|mult_3~124 ;
wire \fp_functions_0|mult_3~125 ;
wire \fp_functions_0|mult_3~126 ;
wire \fp_functions_0|mult_3~127 ;
wire \fp_functions_0|mult_3~128 ;
wire \fp_functions_0|mult_3~129 ;
wire \fp_functions_0|mult_3~130 ;
wire \fp_functions_0|mult_3~131 ;
wire \fp_functions_0|mult_3~132 ;
wire \fp_functions_0|mult_3~133 ;
wire \fp_functions_0|mult_3~134 ;
wire \fp_functions_0|mult_3~135 ;
wire \fp_functions_0|mult_3~136 ;
wire \fp_functions_0|mult_3~137 ;
wire \fp_functions_0|mult_3~138 ;
wire \fp_functions_0|mult_3~139 ;
wire \fp_functions_0|mult_3~140 ;
wire \fp_functions_0|mult_3~141 ;
wire \fp_functions_0|mult_3~142 ;
wire \fp_functions_0|mult_3~143 ;
wire \fp_functions_0|mult_3~144 ;
wire \fp_functions_0|mult_3~145 ;
wire \fp_functions_0|mult_3~146 ;
wire \fp_functions_0|mult_3~147 ;
wire \fp_functions_0|mult_3~148 ;
wire \fp_functions_0|mult_3~149 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_wire[11] ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11~PORTBDATAOUT1 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11~PORTBDATAOUT2 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11~PORTBDATAOUT3 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11~PORTBDATAOUT4 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11~PORTBDATAOUT5 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11~PORTBDATAOUT6 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11~PORTBDATAOUT7 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11~PORTBDATAOUT8 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11~PORTBDATAOUT9 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11~PORTBDATAOUT10 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11~PORTBDATAOUT11 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11~PORTBDATAOUT12 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11~PORTBDATAOUT13 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11~PORTBDATAOUT14 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11~PORTBDATAOUT15 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11~PORTBDATAOUT16 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11~PORTBDATAOUT17 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11~PORTBDATAOUT18 ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11~PORTBDATAOUT19 ;
wire \fp_functions_0|add_7~38_cout ;
wire \fp_functions_0|add_8~38_cout ;
wire \fp_functions_0|add_4~5_sumout ;
wire \fp_functions_0|add_4~6 ;
wire \fp_functions_0|add_4~9_sumout ;
wire \fp_functions_0|add_4~10 ;
wire \fp_functions_0|add_4~13_sumout ;
wire \fp_functions_0|add_4~14 ;
wire \fp_functions_0|add_4~17_sumout ;
wire \fp_functions_0|add_4~18 ;
wire \fp_functions_0|add_4~21_sumout ;
wire \fp_functions_0|add_4~22 ;
wire \fp_functions_0|add_4~25_sumout ;
wire \fp_functions_0|add_4~26 ;
wire \fp_functions_0|add_4~29_sumout ;
wire \fp_functions_0|add_4~30 ;
wire \fp_functions_0|add_4~33_sumout ;
wire \fp_functions_0|add_4~34 ;
wire \fp_functions_0|add_4~37_sumout ;
wire \fp_functions_0|add_4~38 ;
wire \fp_functions_0|add_4~41_sumout ;
wire \fp_functions_0|add_4~42 ;
wire \fp_functions_0|add_7~42_cout ;
wire \fp_functions_0|add_8~42_cout ;
wire \fp_functions_0|add_7~46_cout ;
wire \fp_functions_0|add_8~46_cout ;
wire \fp_functions_0|add_4~45_sumout ;
wire \fp_functions_0|add_7~50_cout ;
wire \fp_functions_0|add_8~50_cout ;
wire \fp_functions_0|add_7~54_cout ;
wire \fp_functions_0|add_8~54_cout ;
wire \fp_functions_0|add_7~58_cout ;
wire \fp_functions_0|add_8~58_cout ;
wire \fp_functions_0|redist10|delay_signals[0][0]~q ;
wire \fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ;
wire \fp_functions_0|ExcROvfAndInReg_uid84_fpMulTest_delay|delay_signals[0][0]~q ;
wire \fp_functions_0|excYRAndExcXI_uid83_fpMulTest_delay|delay_signals[0][0]~q ;
wire \fp_functions_0|excXRAndExcYI_uid82_fpMulTest_delay|delay_signals[0][0]~q ;
wire \fp_functions_0|excXIAndExcYI_uid81_fpMulTest_delay|delay_signals[0][0]~q ;
wire \fp_functions_0|i6400~combout ;
wire \fp_functions_0|excZC3_uid79_fpMulTest_delay|delay_signals[0][0]~q ;
wire \fp_functions_0|excYZAndExcXR_uid78_fpMulTest_delay|delay_signals[0][0]~q ;
wire \fp_functions_0|excXZAndExcYR_uid77_fpMulTest_delay|delay_signals[0][0]~q ;
wire \fp_functions_0|excXZAndExcYZ_uid76_fpMulTest_delay|delay_signals[0][0]~q ;
wire \fp_functions_0|i6475~combout ;
wire \fp_functions_0|Mux_64~0_combout ;
wire \fp_functions_0|redist10|delay_signals[0][1]~q ;
wire \fp_functions_0|Mux_63~0_combout ;
wire \fp_functions_0|redist10|delay_signals[0][2]~q ;
wire \fp_functions_0|Mux_62~0_combout ;
wire \fp_functions_0|redist10|delay_signals[0][3]~q ;
wire \fp_functions_0|Mux_61~0_combout ;
wire \fp_functions_0|redist10|delay_signals[0][4]~q ;
wire \fp_functions_0|Mux_60~0_combout ;
wire \fp_functions_0|redist10|delay_signals[0][5]~q ;
wire \fp_functions_0|Mux_59~0_combout ;
wire \fp_functions_0|redist10|delay_signals[0][6]~q ;
wire \fp_functions_0|Mux_58~0_combout ;
wire \fp_functions_0|redist10|delay_signals[0][7]~q ;
wire \fp_functions_0|Mux_57~0_combout ;
wire \fp_functions_0|redist10|delay_signals[0][8]~q ;
wire \fp_functions_0|Mux_56~0_combout ;
wire \fp_functions_0|redist10|delay_signals[0][9]~q ;
wire \fp_functions_0|Mux_55~0_combout ;
wire \fp_functions_0|redist10|delay_signals[0][10]~q ;
wire \fp_functions_0|Mux_54~0_combout ;
wire \fp_functions_0|redist10|delay_signals[0][11]~q ;
wire \fp_functions_0|Mux_53~0_combout ;
wire \fp_functions_0|redist10|delay_signals[0][12]~q ;
wire \fp_functions_0|Mux_52~0_combout ;
wire \fp_functions_0|redist10|delay_signals[0][13]~q ;
wire \fp_functions_0|Mux_51~0_combout ;
wire \fp_functions_0|redist10|delay_signals[0][14]~q ;
wire \fp_functions_0|Mux_50~0_combout ;
wire \fp_functions_0|redist10|delay_signals[0][15]~q ;
wire \fp_functions_0|Mux_49~0_combout ;
wire \fp_functions_0|redist10|delay_signals[0][16]~q ;
wire \fp_functions_0|Mux_48~0_combout ;
wire \fp_functions_0|redist10|delay_signals[0][17]~q ;
wire \fp_functions_0|Mux_47~0_combout ;
wire \fp_functions_0|redist10|delay_signals[0][18]~q ;
wire \fp_functions_0|Mux_46~0_combout ;
wire \fp_functions_0|redist10|delay_signals[0][19]~q ;
wire \fp_functions_0|Mux_45~0_combout ;
wire \fp_functions_0|redist10|delay_signals[0][20]~q ;
wire \fp_functions_0|Mux_44~0_combout ;
wire \fp_functions_0|redist10|delay_signals[0][21]~q ;
wire \fp_functions_0|Mux_43~0_combout ;
wire \fp_functions_0|redist10|delay_signals[0][22]~q ;
wire \fp_functions_0|Mux_42~0_combout ;
wire \fp_functions_0|redist10|delay_signals[0][23]~q ;
wire \fp_functions_0|Mux_41~0_combout ;
wire \fp_functions_0|redist10|delay_signals[0][24]~q ;
wire \fp_functions_0|Mux_40~0_combout ;
wire \fp_functions_0|redist10|delay_signals[0][25]~q ;
wire \fp_functions_0|Mux_39~0_combout ;
wire \fp_functions_0|redist10|delay_signals[0][26]~q ;
wire \fp_functions_0|Mux_38~0_combout ;
wire \fp_functions_0|redist10|delay_signals[0][27]~q ;
wire \fp_functions_0|Mux_37~0_combout ;
wire \fp_functions_0|redist10|delay_signals[0][28]~q ;
wire \fp_functions_0|Mux_36~0_combout ;
wire \fp_functions_0|redist10|delay_signals[0][29]~q ;
wire \fp_functions_0|Mux_35~0_combout ;
wire \fp_functions_0|redist10|delay_signals[0][30]~q ;
wire \fp_functions_0|Mux_34~0_combout ;
wire \fp_functions_0|redist10|delay_signals[0][31]~q ;
wire \fp_functions_0|Mux_33~0_combout ;
wire \fp_functions_0|redist10|delay_signals[0][32]~q ;
wire \fp_functions_0|Mux_32~0_combout ;
wire \fp_functions_0|redist10|delay_signals[0][33]~q ;
wire \fp_functions_0|Mux_31~0_combout ;
wire \fp_functions_0|redist10|delay_signals[0][34]~q ;
wire \fp_functions_0|Mux_30~0_combout ;
wire \fp_functions_0|redist10|delay_signals[0][35]~q ;
wire \fp_functions_0|Mux_29~0_combout ;
wire \fp_functions_0|redist10|delay_signals[0][36]~q ;
wire \fp_functions_0|Mux_28~0_combout ;
wire \fp_functions_0|redist10|delay_signals[0][37]~q ;
wire \fp_functions_0|Mux_27~0_combout ;
wire \fp_functions_0|redist10|delay_signals[0][38]~q ;
wire \fp_functions_0|Mux_26~0_combout ;
wire \fp_functions_0|redist10|delay_signals[0][39]~q ;
wire \fp_functions_0|Mux_25~0_combout ;
wire \fp_functions_0|redist10|delay_signals[0][40]~q ;
wire \fp_functions_0|Mux_24~0_combout ;
wire \fp_functions_0|redist10|delay_signals[0][41]~q ;
wire \fp_functions_0|Mux_23~0_combout ;
wire \fp_functions_0|redist10|delay_signals[0][42]~q ;
wire \fp_functions_0|Mux_22~0_combout ;
wire \fp_functions_0|redist10|delay_signals[0][43]~q ;
wire \fp_functions_0|Mux_21~0_combout ;
wire \fp_functions_0|redist10|delay_signals[0][44]~q ;
wire \fp_functions_0|Mux_20~0_combout ;
wire \fp_functions_0|redist10|delay_signals[0][45]~q ;
wire \fp_functions_0|Mux_19~0_combout ;
wire \fp_functions_0|redist10|delay_signals[0][46]~q ;
wire \fp_functions_0|Mux_18~0_combout ;
wire \fp_functions_0|redist10|delay_signals[0][47]~q ;
wire \fp_functions_0|Mux_17~0_combout ;
wire \fp_functions_0|redist10|delay_signals[0][48]~q ;
wire \fp_functions_0|Mux_16~0_combout ;
wire \fp_functions_0|redist10|delay_signals[0][49]~q ;
wire \fp_functions_0|Mux_15~0_combout ;
wire \fp_functions_0|redist10|delay_signals[0][50]~q ;
wire \fp_functions_0|Mux_14~0_combout ;
wire \fp_functions_0|redist10|delay_signals[0][51]~q ;
wire \fp_functions_0|Mux_13~0_combout ;
wire \fp_functions_0|redist8|delay_signals[0][0]~q ;
wire \fp_functions_0|Mux_12~0_combout ;
wire \fp_functions_0|redist8|delay_signals[0][1]~q ;
wire \fp_functions_0|Mux_12~1_combout ;
wire \fp_functions_0|redist8|delay_signals[0][2]~q ;
wire \fp_functions_0|Mux_12~2_combout ;
wire \fp_functions_0|redist8|delay_signals[0][3]~q ;
wire \fp_functions_0|Mux_12~3_combout ;
wire \fp_functions_0|redist8|delay_signals[0][4]~q ;
wire \fp_functions_0|Mux_12~4_combout ;
wire \fp_functions_0|redist8|delay_signals[0][5]~q ;
wire \fp_functions_0|Mux_12~5_combout ;
wire \fp_functions_0|redist8|delay_signals[0][6]~q ;
wire \fp_functions_0|Mux_12~6_combout ;
wire \fp_functions_0|redist8|delay_signals[0][7]~q ;
wire \fp_functions_0|Mux_12~7_combout ;
wire \fp_functions_0|redist8|delay_signals[0][8]~q ;
wire \fp_functions_0|Mux_12~8_combout ;
wire \fp_functions_0|redist8|delay_signals[0][9]~q ;
wire \fp_functions_0|Mux_12~9_combout ;
wire \fp_functions_0|redist8|delay_signals[0][10]~q ;
wire \fp_functions_0|Mux_12~10_combout ;
wire \fp_functions_0|redist14|delay_signals[0][0]~q ;
wire \fp_functions_0|i1071~combout ;
wire \fp_functions_0|redist10|delay_signals[1][0]~q ;
wire \fp_functions_0|redist18|delay_signals[0][0]~q ;
wire \fp_functions_0|redist17|delay_signals[0][0]~q ;
wire \fp_functions_0|redist20|delay_signals[0][0]~q ;
wire \fp_functions_0|redist21|delay_signals[0][0]~q ;
wire \fp_functions_0|redist16|delay_signals[0][0]~q ;
wire \fp_functions_0|redist19|delay_signals[0][0]~q ;
wire \fp_functions_0|i933~0_combout ;
wire \fp_functions_0|i6384~combout ;
wire \fp_functions_0|i6387~0_combout ;
wire \fp_functions_0|i6390~0_combout ;
wire \fp_functions_0|i6393~0_combout ;
wire \fp_functions_0|i6459~combout ;
wire \fp_functions_0|i6462~0_combout ;
wire \fp_functions_0|i6465~0_combout ;
wire \fp_functions_0|i6468~combout ;
wire \fp_functions_0|redist10|delay_signals[1][1]~q ;
wire \fp_functions_0|redist10|delay_signals[1][2]~q ;
wire \fp_functions_0|redist10|delay_signals[1][3]~q ;
wire \fp_functions_0|redist10|delay_signals[1][4]~q ;
wire \fp_functions_0|redist10|delay_signals[1][5]~q ;
wire \fp_functions_0|redist10|delay_signals[1][6]~q ;
wire \fp_functions_0|redist10|delay_signals[1][7]~q ;
wire \fp_functions_0|redist10|delay_signals[1][8]~q ;
wire \fp_functions_0|redist10|delay_signals[1][9]~q ;
wire \fp_functions_0|redist10|delay_signals[1][10]~q ;
wire \fp_functions_0|redist10|delay_signals[1][11]~q ;
wire \fp_functions_0|redist10|delay_signals[1][12]~q ;
wire \fp_functions_0|redist10|delay_signals[1][13]~q ;
wire \fp_functions_0|redist10|delay_signals[1][14]~q ;
wire \fp_functions_0|redist10|delay_signals[1][15]~q ;
wire \fp_functions_0|redist10|delay_signals[1][16]~q ;
wire \fp_functions_0|redist10|delay_signals[1][17]~q ;
wire \fp_functions_0|redist10|delay_signals[1][18]~q ;
wire \fp_functions_0|redist10|delay_signals[1][19]~q ;
wire \fp_functions_0|redist10|delay_signals[1][20]~q ;
wire \fp_functions_0|redist10|delay_signals[1][21]~q ;
wire \fp_functions_0|redist10|delay_signals[1][22]~q ;
wire \fp_functions_0|redist10|delay_signals[1][23]~q ;
wire \fp_functions_0|redist10|delay_signals[1][24]~q ;
wire \fp_functions_0|redist10|delay_signals[1][25]~q ;
wire \fp_functions_0|redist10|delay_signals[1][26]~q ;
wire \fp_functions_0|redist10|delay_signals[1][27]~q ;
wire \fp_functions_0|redist10|delay_signals[1][28]~q ;
wire \fp_functions_0|redist10|delay_signals[1][29]~q ;
wire \fp_functions_0|redist10|delay_signals[1][30]~q ;
wire \fp_functions_0|redist10|delay_signals[1][31]~q ;
wire \fp_functions_0|redist10|delay_signals[1][32]~q ;
wire \fp_functions_0|redist10|delay_signals[1][33]~q ;
wire \fp_functions_0|redist10|delay_signals[1][34]~q ;
wire \fp_functions_0|redist10|delay_signals[1][35]~q ;
wire \fp_functions_0|redist10|delay_signals[1][36]~q ;
wire \fp_functions_0|redist10|delay_signals[1][37]~q ;
wire \fp_functions_0|redist10|delay_signals[1][38]~q ;
wire \fp_functions_0|redist10|delay_signals[1][39]~q ;
wire \fp_functions_0|redist10|delay_signals[1][40]~q ;
wire \fp_functions_0|redist10|delay_signals[1][41]~q ;
wire \fp_functions_0|redist10|delay_signals[1][42]~q ;
wire \fp_functions_0|redist10|delay_signals[1][43]~q ;
wire \fp_functions_0|redist10|delay_signals[1][44]~q ;
wire \fp_functions_0|redist10|delay_signals[1][45]~q ;
wire \fp_functions_0|redist10|delay_signals[1][46]~q ;
wire \fp_functions_0|redist10|delay_signals[1][47]~q ;
wire \fp_functions_0|redist10|delay_signals[1][48]~q ;
wire \fp_functions_0|redist10|delay_signals[1][49]~q ;
wire \fp_functions_0|redist10|delay_signals[1][50]~q ;
wire \fp_functions_0|redist10|delay_signals[1][51]~q ;
wire \fp_functions_0|redist9|delay_signals[0][0]~q ;
wire \fp_functions_0|redist9|delay_signals[0][1]~q ;
wire \fp_functions_0|redist9|delay_signals[0][2]~q ;
wire \fp_functions_0|redist9|delay_signals[0][3]~q ;
wire \fp_functions_0|redist9|delay_signals[0][4]~q ;
wire \fp_functions_0|redist9|delay_signals[0][5]~q ;
wire \fp_functions_0|redist9|delay_signals[0][6]~q ;
wire \fp_functions_0|redist9|delay_signals[0][7]~q ;
wire \fp_functions_0|redist9|delay_signals[0][8]~q ;
wire \fp_functions_0|redist9|delay_signals[0][9]~q ;
wire \fp_functions_0|redist9|delay_signals[0][10]~q ;
wire \fp_functions_0|redist14|delay_signals[1][0]~q ;
wire \fp_functions_0|redist18|delay_signals[1][0]~q ;
wire \fp_functions_0|redist17|delay_signals[1][0]~q ;
wire \fp_functions_0|redist20|delay_signals[1][0]~q ;
wire \fp_functions_0|redist21|delay_signals[1][0]~q ;
wire \fp_functions_0|redist16|delay_signals[1][0]~q ;
wire \fp_functions_0|redist19|delay_signals[1][0]~q ;
wire \fp_functions_0|redist9|delay_signals[0][14]~q ;
wire \fp_functions_0|redist14|delay_signals[2][0]~q ;
wire \fp_functions_0|redist11|delay_signals[0][1]~q ;
wire \fp_functions_0|redist18|delay_signals[2][0]~q ;
wire \fp_functions_0|redist17|delay_signals[2][0]~q ;
wire \fp_functions_0|redist20|delay_signals[2][0]~q ;
wire \fp_functions_0|redist21|delay_signals[2][0]~q ;
wire \fp_functions_0|redist16|delay_signals[2][0]~q ;
wire \fp_functions_0|redist19|delay_signals[2][0]~q ;
wire \fp_functions_0|redist11|delay_signals[0][2]~q ;
wire \fp_functions_0|redist11|delay_signals[0][3]~q ;
wire \fp_functions_0|redist11|delay_signals[0][4]~q ;
wire \fp_functions_0|redist11|delay_signals[0][5]~q ;
wire \fp_functions_0|redist11|delay_signals[0][6]~q ;
wire \fp_functions_0|redist11|delay_signals[0][7]~q ;
wire \fp_functions_0|redist11|delay_signals[0][8]~q ;
wire \fp_functions_0|redist11|delay_signals[0][9]~q ;
wire \fp_functions_0|redist11|delay_signals[0][10]~q ;
wire \fp_functions_0|redist11|delay_signals[0][11]~q ;
wire \fp_functions_0|redist11|delay_signals[0][12]~q ;
wire \fp_functions_0|redist11|delay_signals[0][13]~q ;
wire \fp_functions_0|redist11|delay_signals[0][14]~q ;
wire \fp_functions_0|redist11|delay_signals[0][15]~q ;
wire \fp_functions_0|redist11|delay_signals[0][16]~q ;
wire \fp_functions_0|redist11|delay_signals[0][17]~q ;
wire \fp_functions_0|redist11|delay_signals[0][18]~q ;
wire \fp_functions_0|redist11|delay_signals[0][19]~q ;
wire \fp_functions_0|redist11|delay_signals[0][20]~q ;
wire \fp_functions_0|redist11|delay_signals[0][21]~q ;
wire \fp_functions_0|redist11|delay_signals[0][22]~q ;
wire \fp_functions_0|redist11|delay_signals[0][23]~q ;
wire \fp_functions_0|redist11|delay_signals[0][24]~q ;
wire \fp_functions_0|redist11|delay_signals[0][25]~q ;
wire \fp_functions_0|redist11|delay_signals[0][26]~q ;
wire \fp_functions_0|redist11|delay_signals[0][27]~q ;
wire \fp_functions_0|redist11|delay_signals[0][28]~q ;
wire \fp_functions_0|redist11|delay_signals[0][29]~q ;
wire \fp_functions_0|redist11|delay_signals[0][30]~q ;
wire \fp_functions_0|redist11|delay_signals[0][31]~q ;
wire \fp_functions_0|redist11|delay_signals[0][32]~q ;
wire \fp_functions_0|redist11|delay_signals[0][33]~q ;
wire \fp_functions_0|redist11|delay_signals[0][34]~q ;
wire \fp_functions_0|redist11|delay_signals[0][35]~q ;
wire \fp_functions_0|redist11|delay_signals[0][36]~q ;
wire \fp_functions_0|redist11|delay_signals[0][37]~q ;
wire \fp_functions_0|redist11|delay_signals[0][38]~q ;
wire \fp_functions_0|redist11|delay_signals[0][39]~q ;
wire \fp_functions_0|redist11|delay_signals[0][40]~q ;
wire \fp_functions_0|redist11|delay_signals[0][41]~q ;
wire \fp_functions_0|redist11|delay_signals[0][42]~q ;
wire \fp_functions_0|redist11|delay_signals[0][43]~q ;
wire \fp_functions_0|redist11|delay_signals[0][44]~q ;
wire \fp_functions_0|redist11|delay_signals[0][45]~q ;
wire \fp_functions_0|redist11|delay_signals[0][46]~q ;
wire \fp_functions_0|redist11|delay_signals[0][47]~q ;
wire \fp_functions_0|redist11|delay_signals[0][48]~q ;
wire \fp_functions_0|redist11|delay_signals[0][49]~q ;
wire \fp_functions_0|redist11|delay_signals[0][50]~q ;
wire \fp_functions_0|redist11|delay_signals[0][51]~q ;
wire \fp_functions_0|redist11|delay_signals[0][52]~q ;
wire \fp_functions_0|redist11|delay_signals[0][53]~q ;
wire \fp_functions_0|redist13|delay_signals[0][0]~q ;
wire \fp_functions_0|redist11|delay_signals[0][54]~q ;
wire \fp_functions_0|redist11|delay_signals[0][55]~q ;
wire \fp_functions_0|redist11|delay_signals[0][56]~q ;
wire \fp_functions_0|redist11|delay_signals[0][57]~q ;
wire \fp_functions_0|redist11|delay_signals[0][58]~q ;
wire \fp_functions_0|redist11|delay_signals[0][59]~q ;
wire \fp_functions_0|redist11|delay_signals[0][60]~q ;
wire \fp_functions_0|redist11|delay_signals[0][61]~q ;
wire \fp_functions_0|redist11|delay_signals[0][62]~q ;
wire \fp_functions_0|redist11|delay_signals[0][63]~q ;
wire \fp_functions_0|redist14|delay_signals[3][0]~q ;
wire \fp_functions_0|redist11|delay_signals[0][0]~q ;
wire \fp_functions_0|roundBit_uid65_fpMulTest_delay|delay_signals[0][0]~q ;
wire \fp_functions_0|redist18|delay_signals[3][0]~q ;
wire \fp_functions_0|redist17|delay_signals[3][0]~q ;
wire \fp_functions_0|redist20|delay_signals[3][0]~q ;
wire \fp_functions_0|redist21|delay_signals[3][0]~q ;
wire \fp_functions_0|redist16|delay_signals[3][0]~q ;
wire \fp_functions_0|redist19|delay_signals[3][0]~q ;
wire \fp_functions_0|redist11|delay_signals[0][66]~q ;
wire \fp_functions_0|redist9|delay_signals[0][13]~q ;
wire \fp_functions_0|redist15_outputreg|delay_signals[0][0]~q ;
wire \fp_functions_0|redist13|delay_signals[1][0]~q ;
wire \fp_functions_0|redist14|delay_signals[4][0]~q ;
wire \fp_functions_0|redist1|delay_signals[0][52]~q ;
wire \fp_functions_0|redist1|delay_signals[0][53]~q ;
wire \fp_functions_0|redist1|delay_signals[0][105]~q ;
wire \fp_functions_0|redist12|delay_signals[0][48]~q ;
wire \fp_functions_0|redist12|delay_signals[0][49]~q ;
wire \fp_functions_0|redist12|delay_signals[0][50]~q ;
wire \fp_functions_0|redist12|delay_signals[0][51]~q ;
wire \fp_functions_0|reduce_nor_7~0_combout ;
wire \fp_functions_0|redist12|delay_signals[0][41]~q ;
wire \fp_functions_0|redist12|delay_signals[0][46]~q ;
wire \fp_functions_0|redist12|delay_signals[0][47]~q ;
wire \fp_functions_0|redist12|delay_signals[0][42]~q ;
wire \fp_functions_0|redist12|delay_signals[0][43]~q ;
wire \fp_functions_0|redist12|delay_signals[0][44]~q ;
wire \fp_functions_0|redist12|delay_signals[0][45]~q ;
wire \fp_functions_0|reduce_nor_7~1_combout ;
wire \fp_functions_0|redist12|delay_signals[0][36]~q ;
wire \fp_functions_0|redist12|delay_signals[0][37]~q ;
wire \fp_functions_0|redist12|delay_signals[0][38]~q ;
wire \fp_functions_0|redist12|delay_signals[0][39]~q ;
wire \fp_functions_0|redist12|delay_signals[0][40]~q ;
wire \fp_functions_0|reduce_nor_7~2_combout ;
wire \fp_functions_0|reduce_nor_7~3_combout ;
wire \fp_functions_0|redist12|delay_signals[0][29]~q ;
wire \fp_functions_0|redist12|delay_signals[0][35]~q ;
wire \fp_functions_0|redist12|delay_signals[0][24]~q ;
wire \fp_functions_0|redist12|delay_signals[0][25]~q ;
wire \fp_functions_0|redist12|delay_signals[0][26]~q ;
wire \fp_functions_0|redist12|delay_signals[0][27]~q ;
wire \fp_functions_0|redist12|delay_signals[0][28]~q ;
wire \fp_functions_0|reduce_nor_7~4_combout ;
wire \fp_functions_0|redist12|delay_signals[0][30]~q ;
wire \fp_functions_0|redist12|delay_signals[0][31]~q ;
wire \fp_functions_0|redist12|delay_signals[0][32]~q ;
wire \fp_functions_0|redist12|delay_signals[0][33]~q ;
wire \fp_functions_0|redist12|delay_signals[0][34]~q ;
wire \fp_functions_0|reduce_nor_7~5_combout ;
wire \fp_functions_0|redist12|delay_signals[0][17]~q ;
wire \fp_functions_0|redist12|delay_signals[0][23]~q ;
wire \fp_functions_0|redist12|delay_signals[0][12]~q ;
wire \fp_functions_0|redist12|delay_signals[0][13]~q ;
wire \fp_functions_0|redist12|delay_signals[0][14]~q ;
wire \fp_functions_0|redist12|delay_signals[0][15]~q ;
wire \fp_functions_0|redist12|delay_signals[0][16]~q ;
wire \fp_functions_0|reduce_nor_7~6_combout ;
wire \fp_functions_0|redist12|delay_signals[0][18]~q ;
wire \fp_functions_0|redist12|delay_signals[0][19]~q ;
wire \fp_functions_0|redist12|delay_signals[0][20]~q ;
wire \fp_functions_0|redist12|delay_signals[0][21]~q ;
wire \fp_functions_0|redist12|delay_signals[0][22]~q ;
wire \fp_functions_0|reduce_nor_7~7_combout ;
wire \fp_functions_0|redist12|delay_signals[0][5]~q ;
wire \fp_functions_0|redist12|delay_signals[0][10]~q ;
wire \fp_functions_0|redist12|delay_signals[0][11]~q ;
wire \fp_functions_0|redist12|delay_signals[0][6]~q ;
wire \fp_functions_0|redist12|delay_signals[0][7]~q ;
wire \fp_functions_0|redist12|delay_signals[0][8]~q ;
wire \fp_functions_0|redist12|delay_signals[0][9]~q ;
wire \fp_functions_0|reduce_nor_7~8_combout ;
wire \fp_functions_0|redist12|delay_signals[0][0]~q ;
wire \fp_functions_0|redist12|delay_signals[0][1]~q ;
wire \fp_functions_0|redist12|delay_signals[0][2]~q ;
wire \fp_functions_0|redist12|delay_signals[0][3]~q ;
wire \fp_functions_0|redist12|delay_signals[0][4]~q ;
wire \fp_functions_0|reduce_nor_7~9_combout ;
wire \fp_functions_0|reduce_nor_7~10_combout ;
wire \fp_functions_0|reduce_nor_7~combout ;
wire \fp_functions_0|redist18|delay_signals[4][0]~q ;
wire \fp_functions_0|redist17|delay_signals[4][0]~q ;
wire \fp_functions_0|redist20|delay_signals[4][0]~q ;
wire \fp_functions_0|redist21|delay_signals[4][0]~q ;
wire \fp_functions_0|redist16|delay_signals[4][0]~q ;
wire \fp_functions_0|redist19|delay_signals[4][0]~q ;
wire \fp_functions_0|redist9|delay_signals[0][12]~q ;
wire \fp_functions_0|redist1|delay_signals[0][54]~q ;
wire \fp_functions_0|redist1|delay_signals[0][55]~q ;
wire \fp_functions_0|redist1|delay_signals[0][56]~q ;
wire \fp_functions_0|redist1|delay_signals[0][57]~q ;
wire \fp_functions_0|redist1|delay_signals[0][58]~q ;
wire \fp_functions_0|redist1|delay_signals[0][59]~q ;
wire \fp_functions_0|redist1|delay_signals[0][60]~q ;
wire \fp_functions_0|redist1|delay_signals[0][61]~q ;
wire \fp_functions_0|redist1|delay_signals[0][62]~q ;
wire \fp_functions_0|redist1|delay_signals[0][63]~q ;
wire \fp_functions_0|redist1|delay_signals[0][64]~q ;
wire \fp_functions_0|redist1|delay_signals[0][65]~q ;
wire \fp_functions_0|redist1|delay_signals[0][66]~q ;
wire \fp_functions_0|redist1|delay_signals[0][67]~q ;
wire \fp_functions_0|redist1|delay_signals[0][68]~q ;
wire \fp_functions_0|redist1|delay_signals[0][69]~q ;
wire \fp_functions_0|redist1|delay_signals[0][70]~q ;
wire \fp_functions_0|redist1|delay_signals[0][71]~q ;
wire \fp_functions_0|redist1|delay_signals[0][72]~q ;
wire \fp_functions_0|redist1|delay_signals[0][73]~q ;
wire \fp_functions_0|redist1|delay_signals[0][74]~q ;
wire \fp_functions_0|redist1|delay_signals[0][75]~q ;
wire \fp_functions_0|redist1|delay_signals[0][76]~q ;
wire \fp_functions_0|redist1|delay_signals[0][77]~q ;
wire \fp_functions_0|redist1|delay_signals[0][78]~q ;
wire \fp_functions_0|redist1|delay_signals[0][79]~q ;
wire \fp_functions_0|redist1|delay_signals[0][80]~q ;
wire \fp_functions_0|redist1|delay_signals[0][81]~q ;
wire \fp_functions_0|redist1|delay_signals[0][82]~q ;
wire \fp_functions_0|redist1|delay_signals[0][83]~q ;
wire \fp_functions_0|redist1|delay_signals[0][84]~q ;
wire \fp_functions_0|redist1|delay_signals[0][85]~q ;
wire \fp_functions_0|redist1|delay_signals[0][86]~q ;
wire \fp_functions_0|redist1|delay_signals[0][87]~q ;
wire \fp_functions_0|redist1|delay_signals[0][88]~q ;
wire \fp_functions_0|redist1|delay_signals[0][89]~q ;
wire \fp_functions_0|redist1|delay_signals[0][90]~q ;
wire \fp_functions_0|redist1|delay_signals[0][91]~q ;
wire \fp_functions_0|redist1|delay_signals[0][92]~q ;
wire \fp_functions_0|redist1|delay_signals[0][93]~q ;
wire \fp_functions_0|redist1|delay_signals[0][94]~q ;
wire \fp_functions_0|redist1|delay_signals[0][95]~q ;
wire \fp_functions_0|redist1|delay_signals[0][96]~q ;
wire \fp_functions_0|redist1|delay_signals[0][97]~q ;
wire \fp_functions_0|redist1|delay_signals[0][98]~q ;
wire \fp_functions_0|redist1|delay_signals[0][99]~q ;
wire \fp_functions_0|redist1|delay_signals[0][100]~q ;
wire \fp_functions_0|redist1|delay_signals[0][101]~q ;
wire \fp_functions_0|redist1|delay_signals[0][102]~q ;
wire \fp_functions_0|redist1|delay_signals[0][103]~q ;
wire \fp_functions_0|redist1|delay_signals[0][104]~q ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[0]~q ;
wire \fp_functions_0|redist15_outputreg|delay_signals[0][1]~q ;
wire \fp_functions_0|redist15_outputreg|delay_signals[0][2]~q ;
wire \fp_functions_0|redist15_outputreg|delay_signals[0][3]~q ;
wire \fp_functions_0|redist15_outputreg|delay_signals[0][4]~q ;
wire \fp_functions_0|redist15_outputreg|delay_signals[0][5]~q ;
wire \fp_functions_0|redist15_outputreg|delay_signals[0][6]~q ;
wire \fp_functions_0|redist15_outputreg|delay_signals[0][7]~q ;
wire \fp_functions_0|redist15_outputreg|delay_signals[0][8]~q ;
wire \fp_functions_0|redist15_outputreg|delay_signals[0][9]~q ;
wire \fp_functions_0|redist15_outputreg|delay_signals[0][10]~q ;
wire \fp_functions_0|redist14|delay_signals[5][0]~q ;
wire \fp_functions_0|redist1|delay_signals[0][51]~q ;
wire \fp_functions_0|redist1|delay_signals[0][48]~q ;
wire \fp_functions_0|redist1|delay_signals[0][49]~q ;
wire \fp_functions_0|redist1|delay_signals[0][50]~q ;
wire \fp_functions_0|i5343~0_combout ;
wire \fp_functions_0|redist1|delay_signals[0][41]~q ;
wire \fp_functions_0|redist1|delay_signals[0][46]~q ;
wire \fp_functions_0|redist1|delay_signals[0][47]~q ;
wire \fp_functions_0|redist1|delay_signals[0][42]~q ;
wire \fp_functions_0|redist1|delay_signals[0][43]~q ;
wire \fp_functions_0|redist1|delay_signals[0][44]~q ;
wire \fp_functions_0|redist1|delay_signals[0][45]~q ;
wire \fp_functions_0|redist1|delay_signals[0][36]~q ;
wire \fp_functions_0|redist1|delay_signals[0][37]~q ;
wire \fp_functions_0|redist1|delay_signals[0][38]~q ;
wire \fp_functions_0|redist1|delay_signals[0][39]~q ;
wire \fp_functions_0|redist1|delay_signals[0][40]~q ;
wire \fp_functions_0|redist1|delay_signals[0][29]~q ;
wire \fp_functions_0|redist1|delay_signals[0][35]~q ;
wire \fp_functions_0|redist1|delay_signals[0][24]~q ;
wire \fp_functions_0|redist1|delay_signals[0][25]~q ;
wire \fp_functions_0|redist1|delay_signals[0][26]~q ;
wire \fp_functions_0|redist1|delay_signals[0][27]~q ;
wire \fp_functions_0|redist1|delay_signals[0][28]~q ;
wire \fp_functions_0|redist1|delay_signals[0][30]~q ;
wire \fp_functions_0|redist1|delay_signals[0][31]~q ;
wire \fp_functions_0|redist1|delay_signals[0][32]~q ;
wire \fp_functions_0|redist1|delay_signals[0][33]~q ;
wire \fp_functions_0|redist1|delay_signals[0][34]~q ;
wire \fp_functions_0|redist1|delay_signals[0][17]~q ;
wire \fp_functions_0|redist1|delay_signals[0][23]~q ;
wire \fp_functions_0|redist1|delay_signals[0][12]~q ;
wire \fp_functions_0|redist1|delay_signals[0][13]~q ;
wire \fp_functions_0|redist1|delay_signals[0][14]~q ;
wire \fp_functions_0|redist1|delay_signals[0][15]~q ;
wire \fp_functions_0|redist1|delay_signals[0][16]~q ;
wire \fp_functions_0|redist1|delay_signals[0][18]~q ;
wire \fp_functions_0|redist1|delay_signals[0][19]~q ;
wire \fp_functions_0|redist1|delay_signals[0][20]~q ;
wire \fp_functions_0|redist1|delay_signals[0][21]~q ;
wire \fp_functions_0|redist1|delay_signals[0][22]~q ;
wire \fp_functions_0|redist1|delay_signals[0][5]~q ;
wire \fp_functions_0|redist1|delay_signals[0][10]~q ;
wire \fp_functions_0|redist1|delay_signals[0][11]~q ;
wire \fp_functions_0|redist1|delay_signals[0][6]~q ;
wire \fp_functions_0|redist1|delay_signals[0][7]~q ;
wire \fp_functions_0|redist1|delay_signals[0][8]~q ;
wire \fp_functions_0|redist1|delay_signals[0][9]~q ;
wire \fp_functions_0|redist1|delay_signals[0][0]~q ;
wire \fp_functions_0|redist1|delay_signals[0][1]~q ;
wire \fp_functions_0|redist1|delay_signals[0][2]~q ;
wire \fp_functions_0|redist1|delay_signals[0][3]~q ;
wire \fp_functions_0|redist1|delay_signals[0][4]~q ;
wire \fp_functions_0|redist18|delay_signals[5][0]~q ;
wire \fp_functions_0|redist17|delay_signals[5][0]~q ;
wire \fp_functions_0|redist20|delay_signals[5][0]~q ;
wire \fp_functions_0|redist21|delay_signals[5][0]~q ;
wire \fp_functions_0|redist16|delay_signals[5][0]~q ;
wire \fp_functions_0|redist19|delay_signals[5][0]~q ;
wire \fp_functions_0|redist11|delay_signals[0][65]~q ;
wire \fp_functions_0|redist9|delay_signals[0][11]~q ;
wire \fp_functions_0|redist15_sticky_ena_q[0]~q ;
wire \fp_functions_0|i5762~combout ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[1]~q ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[2]~q ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[3]~q ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[4]~q ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[5]~q ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[6]~q ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[7]~q ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[8]~q ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[9]~q ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[10]~q ;
wire \fp_functions_0|redist14|delay_signals[6][0]~q ;
wire \fp_functions_0|redist0|delay_signals[0][27]~q ;
wire \fp_functions_0|redist2|delay_signals[0][27]~q ;
wire \fp_functions_0|redist0|delay_signals[0][28]~q ;
wire \fp_functions_0|redist2|delay_signals[0][28]~q ;
wire \fp_functions_0|redist2|delay_signals[0][80]~q ;
wire \fp_functions_0|redist3|delay_signals[0][26]~q ;
wire \fp_functions_0|redist3|delay_signals[0][19]~q ;
wire \fp_functions_0|redist3|delay_signals[0][25]~q ;
wire \fp_functions_0|redist3|delay_signals[0][14]~q ;
wire \fp_functions_0|redist3|delay_signals[0][15]~q ;
wire \fp_functions_0|redist3|delay_signals[0][16]~q ;
wire \fp_functions_0|redist3|delay_signals[0][17]~q ;
wire \fp_functions_0|redist3|delay_signals[0][18]~q ;
wire \fp_functions_0|redist3|delay_signals[0][20]~q ;
wire \fp_functions_0|redist3|delay_signals[0][21]~q ;
wire \fp_functions_0|redist3|delay_signals[0][22]~q ;
wire \fp_functions_0|redist3|delay_signals[0][23]~q ;
wire \fp_functions_0|redist3|delay_signals[0][24]~q ;
wire \fp_functions_0|redist3|delay_signals[0][7]~q ;
wire \fp_functions_0|redist3|delay_signals[0][12]~q ;
wire \fp_functions_0|redist3|delay_signals[0][13]~q ;
wire \fp_functions_0|redist3|delay_signals[0][8]~q ;
wire \fp_functions_0|redist3|delay_signals[0][9]~q ;
wire \fp_functions_0|redist3|delay_signals[0][10]~q ;
wire \fp_functions_0|redist3|delay_signals[0][11]~q ;
wire \fp_functions_0|redist3|delay_signals[0][2]~q ;
wire \fp_functions_0|redist3|delay_signals[0][3]~q ;
wire \fp_functions_0|redist3|delay_signals[0][4]~q ;
wire \fp_functions_0|redist3|delay_signals[0][5]~q ;
wire \fp_functions_0|redist3|delay_signals[0][6]~q ;
wire \fp_functions_0|redist18|delay_signals[6][0]~q ;
wire \fp_functions_0|redist17|delay_signals[6][0]~q ;
wire \fp_functions_0|redist20|delay_signals[6][0]~q ;
wire \fp_functions_0|redist21|delay_signals[6][0]~q ;
wire \fp_functions_0|redist16|delay_signals[6][0]~q ;
wire \fp_functions_0|redist19|delay_signals[6][0]~q ;
wire \fp_functions_0|redist11|delay_signals[0][64]~q ;
wire \fp_functions_0|redist0|delay_signals[0][29]~q ;
wire \fp_functions_0|redist2|delay_signals[0][29]~q ;
wire \fp_functions_0|redist0|delay_signals[0][30]~q ;
wire \fp_functions_0|redist2|delay_signals[0][30]~q ;
wire \fp_functions_0|redist0|delay_signals[0][31]~q ;
wire \fp_functions_0|redist2|delay_signals[0][31]~q ;
wire \fp_functions_0|redist0|delay_signals[0][32]~q ;
wire \fp_functions_0|redist2|delay_signals[0][32]~q ;
wire \fp_functions_0|redist0|delay_signals[0][33]~q ;
wire \fp_functions_0|redist2|delay_signals[0][33]~q ;
wire \fp_functions_0|redist0|delay_signals[0][34]~q ;
wire \fp_functions_0|redist2|delay_signals[0][34]~q ;
wire \fp_functions_0|redist0|delay_signals[0][35]~q ;
wire \fp_functions_0|redist2|delay_signals[0][35]~q ;
wire \fp_functions_0|redist0|delay_signals[0][36]~q ;
wire \fp_functions_0|redist2|delay_signals[0][36]~q ;
wire \fp_functions_0|redist0|delay_signals[0][37]~q ;
wire \fp_functions_0|redist2|delay_signals[0][37]~q ;
wire \fp_functions_0|redist0|delay_signals[0][38]~q ;
wire \fp_functions_0|redist2|delay_signals[0][38]~q ;
wire \fp_functions_0|redist0|delay_signals[0][39]~q ;
wire \fp_functions_0|redist2|delay_signals[0][39]~q ;
wire \fp_functions_0|redist0|delay_signals[0][40]~q ;
wire \fp_functions_0|redist2|delay_signals[0][40]~q ;
wire \fp_functions_0|redist0|delay_signals[0][41]~q ;
wire \fp_functions_0|redist2|delay_signals[0][41]~q ;
wire \fp_functions_0|redist0|delay_signals[0][42]~q ;
wire \fp_functions_0|redist2|delay_signals[0][42]~q ;
wire \fp_functions_0|redist0|delay_signals[0][43]~q ;
wire \fp_functions_0|redist2|delay_signals[0][43]~q ;
wire \fp_functions_0|redist0|delay_signals[0][44]~q ;
wire \fp_functions_0|redist2|delay_signals[0][44]~q ;
wire \fp_functions_0|redist0|delay_signals[0][45]~q ;
wire \fp_functions_0|redist2|delay_signals[0][45]~q ;
wire \fp_functions_0|redist0|delay_signals[0][46]~q ;
wire \fp_functions_0|redist2|delay_signals[0][46]~q ;
wire \fp_functions_0|redist0|delay_signals[0][47]~q ;
wire \fp_functions_0|redist2|delay_signals[0][47]~q ;
wire \fp_functions_0|redist0|delay_signals[0][48]~q ;
wire \fp_functions_0|redist2|delay_signals[0][48]~q ;
wire \fp_functions_0|redist0|delay_signals[0][49]~q ;
wire \fp_functions_0|redist2|delay_signals[0][49]~q ;
wire \fp_functions_0|redist0|delay_signals[0][50]~q ;
wire \fp_functions_0|redist2|delay_signals[0][50]~q ;
wire \fp_functions_0|redist0|delay_signals[0][51]~q ;
wire \fp_functions_0|redist2|delay_signals[0][51]~q ;
wire \fp_functions_0|redist0|delay_signals[0][52]~q ;
wire \fp_functions_0|redist2|delay_signals[0][52]~q ;
wire \fp_functions_0|redist0|delay_signals[0][53]~q ;
wire \fp_functions_0|redist2|delay_signals[0][53]~q ;
wire \fp_functions_0|redist0|delay_signals[0][54]~q ;
wire \fp_functions_0|redist2|delay_signals[0][54]~q ;
wire \fp_functions_0|redist2|delay_signals[0][55]~q ;
wire \fp_functions_0|redist2|delay_signals[0][56]~q ;
wire \fp_functions_0|redist2|delay_signals[0][57]~q ;
wire \fp_functions_0|redist2|delay_signals[0][58]~q ;
wire \fp_functions_0|redist2|delay_signals[0][59]~q ;
wire \fp_functions_0|redist2|delay_signals[0][60]~q ;
wire \fp_functions_0|redist2|delay_signals[0][61]~q ;
wire \fp_functions_0|redist2|delay_signals[0][62]~q ;
wire \fp_functions_0|redist2|delay_signals[0][63]~q ;
wire \fp_functions_0|redist2|delay_signals[0][64]~q ;
wire \fp_functions_0|redist2|delay_signals[0][65]~q ;
wire \fp_functions_0|redist2|delay_signals[0][66]~q ;
wire \fp_functions_0|redist2|delay_signals[0][67]~q ;
wire \fp_functions_0|redist2|delay_signals[0][68]~q ;
wire \fp_functions_0|redist2|delay_signals[0][69]~q ;
wire \fp_functions_0|redist2|delay_signals[0][70]~q ;
wire \fp_functions_0|redist2|delay_signals[0][71]~q ;
wire \fp_functions_0|redist2|delay_signals[0][72]~q ;
wire \fp_functions_0|redist2|delay_signals[0][73]~q ;
wire \fp_functions_0|redist2|delay_signals[0][74]~q ;
wire \fp_functions_0|redist2|delay_signals[0][75]~q ;
wire \fp_functions_0|redist2|delay_signals[0][76]~q ;
wire \fp_functions_0|redist2|delay_signals[0][77]~q ;
wire \fp_functions_0|redist2|delay_signals[0][78]~q ;
wire \fp_functions_0|redist2|delay_signals[0][79]~q ;
wire \fp_functions_0|redist15_wraddr_q[0]~q ;
wire \fp_functions_0|redist15_wraddr_q[1]~q ;
wire \fp_functions_0|redist15_inputreg|delay_signals[0][0]~q ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|rdaddr_reg[0]~q ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|rdaddr_reg[1]~q ;
wire \fp_functions_0|redist15_cmpReg_q[0]~q ;
wire \fp_functions_0|redist15_sticky_ena_q[0]~0_combout ;
wire \fp_functions_0|redist14|delay_signals[7][0]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][27]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][0]~q ;
wire \fp_functions_0|redist0|delay_signals[0][26]~q ;
wire \fp_functions_0|redist2|delay_signals[0][26]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][28]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][1]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][53]~q ;
wire \fp_functions_0|redist0|delay_signals[0][23]~q ;
wire \fp_functions_0|redist2|delay_signals[0][23]~q ;
wire \fp_functions_0|redist0|delay_signals[0][24]~q ;
wire \fp_functions_0|redist2|delay_signals[0][24]~q ;
wire \fp_functions_0|redist0|delay_signals[0][25]~q ;
wire \fp_functions_0|redist2|delay_signals[0][25]~q ;
wire \fp_functions_0|redist0|delay_signals[0][16]~q ;
wire \fp_functions_0|redist2|delay_signals[0][16]~q ;
wire \fp_functions_0|redist0|delay_signals[0][21]~q ;
wire \fp_functions_0|redist2|delay_signals[0][21]~q ;
wire \fp_functions_0|redist0|delay_signals[0][22]~q ;
wire \fp_functions_0|redist2|delay_signals[0][22]~q ;
wire \fp_functions_0|redist0|delay_signals[0][17]~q ;
wire \fp_functions_0|redist2|delay_signals[0][17]~q ;
wire \fp_functions_0|redist0|delay_signals[0][18]~q ;
wire \fp_functions_0|redist2|delay_signals[0][18]~q ;
wire \fp_functions_0|redist0|delay_signals[0][19]~q ;
wire \fp_functions_0|redist2|delay_signals[0][19]~q ;
wire \fp_functions_0|redist0|delay_signals[0][20]~q ;
wire \fp_functions_0|redist2|delay_signals[0][20]~q ;
wire \fp_functions_0|redist0|delay_signals[0][11]~q ;
wire \fp_functions_0|redist2|delay_signals[0][11]~q ;
wire \fp_functions_0|redist0|delay_signals[0][12]~q ;
wire \fp_functions_0|redist2|delay_signals[0][12]~q ;
wire \fp_functions_0|redist0|delay_signals[0][13]~q ;
wire \fp_functions_0|redist2|delay_signals[0][13]~q ;
wire \fp_functions_0|redist0|delay_signals[0][14]~q ;
wire \fp_functions_0|redist2|delay_signals[0][14]~q ;
wire \fp_functions_0|redist0|delay_signals[0][15]~q ;
wire \fp_functions_0|redist2|delay_signals[0][15]~q ;
wire \fp_functions_0|redist0|delay_signals[0][4]~q ;
wire \fp_functions_0|redist2|delay_signals[0][4]~q ;
wire \fp_functions_0|redist0|delay_signals[0][10]~q ;
wire \fp_functions_0|redist2|delay_signals[0][10]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][26]~q ;
wire \fp_functions_0|redist0|delay_signals[0][0]~q ;
wire \fp_functions_0|redist2|delay_signals[0][0]~q ;
wire \fp_functions_0|redist0|delay_signals[0][1]~q ;
wire \fp_functions_0|redist2|delay_signals[0][1]~q ;
wire \fp_functions_0|redist0|delay_signals[0][2]~q ;
wire \fp_functions_0|redist2|delay_signals[0][2]~q ;
wire \fp_functions_0|redist0|delay_signals[0][3]~q ;
wire \fp_functions_0|redist2|delay_signals[0][3]~q ;
wire \fp_functions_0|redist0|delay_signals[0][5]~q ;
wire \fp_functions_0|redist2|delay_signals[0][5]~q ;
wire \fp_functions_0|redist0|delay_signals[0][6]~q ;
wire \fp_functions_0|redist2|delay_signals[0][6]~q ;
wire \fp_functions_0|redist0|delay_signals[0][7]~q ;
wire \fp_functions_0|redist2|delay_signals[0][7]~q ;
wire \fp_functions_0|redist0|delay_signals[0][8]~q ;
wire \fp_functions_0|redist2|delay_signals[0][8]~q ;
wire \fp_functions_0|redist0|delay_signals[0][9]~q ;
wire \fp_functions_0|redist2|delay_signals[0][9]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][19]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][25]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][14]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][15]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][16]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][17]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][18]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][20]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][21]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][22]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][23]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][24]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][7]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][12]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][13]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][8]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][9]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][10]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][11]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][2]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][3]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][4]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][5]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][6]~q ;
wire \fp_functions_0|redist18|delay_signals[7][0]~q ;
wire \fp_functions_0|redist17|delay_signals[7][0]~q ;
wire \fp_functions_0|redist20|delay_signals[7][0]~q ;
wire \fp_functions_0|redist21|delay_signals[7][0]~q ;
wire \fp_functions_0|redist16|delay_signals[7][0]~q ;
wire \fp_functions_0|redist19|delay_signals[7][0]~q ;
wire \fp_functions_0|redist15_outputreg|delay_signals[0][11]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][29]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][2]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][30]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][3]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][31]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][4]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][32]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][5]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][33]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][6]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][34]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][7]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][35]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][8]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][36]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][9]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][37]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][10]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][38]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][11]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][39]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][12]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][40]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][13]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][41]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][14]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][42]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][15]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][43]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][16]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][44]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][17]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][45]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][18]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][46]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][19]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][47]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][20]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][48]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][21]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][49]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][22]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][50]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][23]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][51]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][24]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][52]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][25]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][53]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][26]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][54]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][27]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][28]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][29]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][30]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][31]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][32]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][33]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][34]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][35]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][36]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][37]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][38]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][39]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][40]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][41]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][42]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][43]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][44]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][45]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][46]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][47]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][48]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][49]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][50]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][51]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][52]~q ;
wire \fp_functions_0|redist15_rdcnt_i[0]~q ;
wire \fp_functions_0|i5779~0_combout ;
wire \fp_functions_0|redist15_rdcnt_i[1]~q ;
wire \fp_functions_0|i5779~1_combout ;
wire \fp_functions_0|expSum_uid44_fpMulTest_o[0]~q ;
wire \fp_functions_0|reduce_nor_8~combout ;
wire \fp_functions_0|redist15_inputreg|delay_signals[0][1]~q ;
wire \fp_functions_0|redist15_inputreg|delay_signals[0][2]~q ;
wire \fp_functions_0|redist15_inputreg|delay_signals[0][3]~q ;
wire \fp_functions_0|redist15_inputreg|delay_signals[0][4]~q ;
wire \fp_functions_0|redist15_inputreg|delay_signals[0][5]~q ;
wire \fp_functions_0|redist15_inputreg|delay_signals[0][6]~q ;
wire \fp_functions_0|redist15_inputreg|delay_signals[0][7]~q ;
wire \fp_functions_0|redist15_inputreg|delay_signals[0][8]~q ;
wire \fp_functions_0|redist15_inputreg|delay_signals[0][9]~q ;
wire \fp_functions_0|redist15_inputreg|delay_signals[0][10]~q ;
wire \fp_functions_0|redist14|delay_signals[8][0]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][26]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][53]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][23]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][50]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][24]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][51]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][25]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][52]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][16]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][43]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][21]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][48]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][22]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][49]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][17]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][44]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][18]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][45]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][19]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][46]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][20]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][47]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][11]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][38]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][12]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][39]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][13]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][40]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][14]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][41]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][15]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][42]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][4]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][31]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][10]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][37]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][0]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][27]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][1]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][28]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][2]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][29]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][3]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][30]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][5]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][32]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][6]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][33]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][7]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][34]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][8]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][35]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][9]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][36]~q ;
wire \fp_functions_0|excZ_y_uid29_fpMulTest_delay|delay_signals[0][0]~q ;
wire \fp_functions_0|expXIsMax_uid30_fpMulTest_delay|delay_signals[0][0]~q ;
wire \fp_functions_0|expXIsMax_uid16_fpMulTest_delay|delay_signals[0][0]~q ;
wire \fp_functions_0|excZ_x_uid15_fpMulTest_delay|delay_signals[0][0]~q ;
wire \fp_functions_0|fracXIsZero_uid31_fpMulTest_delay|delay_signals[0][0]~q ;
wire \fp_functions_0|fracXIsZero_uid17_fpMulTest_delay|delay_signals[0][0]~q ;
wire \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[11]~q ;
wire \fp_functions_0|redist15_rdcnt_eq~q ;
wire \fp_functions_0|redist15_rdcnt_i[0]~0_combout ;
wire \fp_functions_0|i5766~0_combout ;
wire \fp_functions_0|expSum_uid44_fpMulTest_o[1]~q ;
wire \fp_functions_0|expSum_uid44_fpMulTest_o[2]~q ;
wire \fp_functions_0|expSum_uid44_fpMulTest_o[3]~q ;
wire \fp_functions_0|expSum_uid44_fpMulTest_o[4]~q ;
wire \fp_functions_0|expSum_uid44_fpMulTest_o[5]~q ;
wire \fp_functions_0|expSum_uid44_fpMulTest_o[6]~q ;
wire \fp_functions_0|expSum_uid44_fpMulTest_o[7]~q ;
wire \fp_functions_0|expSum_uid44_fpMulTest_o[8]~q ;
wire \fp_functions_0|expSum_uid44_fpMulTest_o[9]~q ;
wire \fp_functions_0|expSum_uid44_fpMulTest_o[10]~q ;
wire \fp_functions_0|signR_uid48_fpMulTest_delay|delay_signals[0][0]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][0]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][1]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][2]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][3]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][4]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][5]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][6]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][7]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][8]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][9]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][10]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][11]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][12]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][13]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][14]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][15]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][16]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][17]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][18]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][19]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][20]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][21]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][22]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][23]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][24]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][25]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][26]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][0]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][1]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][2]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][3]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][4]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][5]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][6]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][7]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][8]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][9]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][10]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][11]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][12]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][13]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][14]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][15]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][16]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][17]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][18]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][19]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][20]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][21]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][22]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][23]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][24]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][25]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][26]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][0]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][1]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][2]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][3]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][4]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][5]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][6]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][7]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][8]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][9]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][10]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][11]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][12]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][13]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][14]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][15]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][16]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][17]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][18]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][19]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][20]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][21]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][22]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][23]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][24]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][25]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][26]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][0]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][1]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][2]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][3]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][4]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][5]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][6]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][7]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][8]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][9]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][10]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][11]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][12]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][13]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][14]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][15]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][16]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][17]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][18]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][19]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][20]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][21]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][22]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][23]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][24]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][25]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][26]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][0]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][1]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][2]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][3]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][4]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][5]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][6]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][7]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][8]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][9]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][10]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][11]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][12]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][13]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][14]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][15]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][16]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][17]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][18]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][19]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][20]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][21]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][22]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][23]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][24]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][25]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][26]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][0]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][1]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][2]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][3]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][4]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][5]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][6]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][7]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][8]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][9]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][10]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][11]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][12]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][13]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][14]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][15]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][16]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][17]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][18]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][19]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][20]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][21]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][22]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][23]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][24]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][25]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][26]~q ;
wire \fp_functions_0|reduce_nor_2~0_combout ;
wire \fp_functions_0|reduce_nor_2~1_combout ;
wire \fp_functions_0|reduce_nor_2~combout ;
wire \fp_functions_0|reduce_nor_4~0_combout ;
wire \fp_functions_0|reduce_nor_4~1_combout ;
wire \fp_functions_0|reduce_nor_4~combout ;
wire \fp_functions_0|reduce_nor_1~0_combout ;
wire \fp_functions_0|reduce_nor_1~1_combout ;
wire \fp_functions_0|reduce_nor_1~combout ;
wire \fp_functions_0|reduce_nor_5~0_combout ;
wire \fp_functions_0|reduce_nor_5~1_combout ;
wire \fp_functions_0|reduce_nor_5~combout ;
wire \fp_functions_0|reduce_nor_3~0_combout ;
wire \fp_functions_0|reduce_nor_3~1_combout ;
wire \fp_functions_0|reduce_nor_3~2_combout ;
wire \fp_functions_0|reduce_nor_3~3_combout ;
wire \fp_functions_0|reduce_nor_3~4_combout ;
wire \fp_functions_0|reduce_nor_3~5_combout ;
wire \fp_functions_0|reduce_nor_3~6_combout ;
wire \fp_functions_0|reduce_nor_3~7_combout ;
wire \fp_functions_0|reduce_nor_3~8_combout ;
wire \fp_functions_0|reduce_nor_3~9_combout ;
wire \fp_functions_0|reduce_nor_3~10_combout ;
wire \fp_functions_0|reduce_nor_3~combout ;
wire \fp_functions_0|reduce_nor_0~0_combout ;
wire \fp_functions_0|reduce_nor_0~1_combout ;
wire \fp_functions_0|reduce_nor_0~2_combout ;
wire \fp_functions_0|reduce_nor_0~3_combout ;
wire \fp_functions_0|reduce_nor_0~4_combout ;
wire \fp_functions_0|reduce_nor_0~5_combout ;
wire \fp_functions_0|reduce_nor_0~6_combout ;
wire \fp_functions_0|reduce_nor_0~7_combout ;
wire \fp_functions_0|reduce_nor_0~8_combout ;
wire \fp_functions_0|reduce_nor_0~9_combout ;
wire \fp_functions_0|reduce_nor_0~10_combout ;
wire \fp_functions_0|reduce_nor_0~combout ;
wire \fp_functions_0|reduce_nor_9~combout ;
wire \fp_functions_0|i1068~combout ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][0]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][1]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][2]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][3]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][4]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][5]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][6]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][7]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][8]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][9]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][10]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][11]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][12]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][13]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][14]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][15]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][16]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][17]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][18]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][19]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][20]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][21]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][22]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][23]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][24]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][25]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][26]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][0]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][1]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][2]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][3]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][4]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][5]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][6]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][7]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][8]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][9]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][10]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][11]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][12]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][13]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][14]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][15]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][16]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][17]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][18]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][19]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][20]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][21]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][22]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][23]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][24]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][25]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][26]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][0]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][1]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][2]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][3]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][4]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][5]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][6]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][7]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][8]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][9]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][10]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][11]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][12]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][13]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][14]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][15]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][16]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][17]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][18]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][19]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][20]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][21]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][22]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][23]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][24]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][25]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][26]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][0]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][1]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][2]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][3]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][4]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][5]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][6]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][7]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][8]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][9]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][10]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][11]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][12]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][13]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][14]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][15]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][16]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][17]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][18]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][19]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][20]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][21]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][22]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][23]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][24]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][25]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][26]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][0]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][1]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][2]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][3]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][4]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][5]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][6]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][7]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][8]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][9]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][10]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][11]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][12]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][13]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][14]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][15]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][16]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][17]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][18]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][19]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][20]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][21]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][22]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][23]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][24]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][25]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][26]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][0]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][1]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][2]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][3]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][4]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][5]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][6]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][7]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][8]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][9]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][10]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][11]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][12]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][13]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][14]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][15]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][16]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][17]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][18]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][19]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][20]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][21]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][22]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][23]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][24]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][25]~q ;
wire \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][26]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][0]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][1]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][2]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][3]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][4]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][5]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][6]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][7]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][8]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][9]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][10]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][11]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][12]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][13]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][14]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][15]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][16]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][17]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][18]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][19]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][20]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][21]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][22]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][23]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][24]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][25]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][26]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][0]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][1]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][2]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][3]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][4]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][5]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][6]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][7]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][8]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][9]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][10]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][11]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][12]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][13]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][14]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][15]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][16]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][17]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][18]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][19]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][20]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][21]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][22]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][23]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][24]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][25]~q ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][26]~q ;
wire \fp_functions_0|redist15_inputreg|delay_signals[0][11]~q ;
wire \fp_functions_0|redist6|delay_signals[0][0]~q ;
wire \fp_functions_0|redist6|delay_signals[0][1]~q ;
wire \fp_functions_0|redist6|delay_signals[0][2]~q ;
wire \fp_functions_0|redist6|delay_signals[0][3]~q ;
wire \fp_functions_0|redist6|delay_signals[0][4]~q ;
wire \fp_functions_0|redist6|delay_signals[0][5]~q ;
wire \fp_functions_0|redist6|delay_signals[0][6]~q ;
wire \fp_functions_0|redist6|delay_signals[0][7]~q ;
wire \fp_functions_0|redist6|delay_signals[0][8]~q ;
wire \fp_functions_0|redist6|delay_signals[0][9]~q ;
wire \fp_functions_0|redist6|delay_signals[0][10]~q ;
wire \fp_functions_0|redist6|delay_signals[0][11]~q ;
wire \fp_functions_0|redist6|delay_signals[0][12]~q ;
wire \fp_functions_0|redist6|delay_signals[0][13]~q ;
wire \fp_functions_0|redist6|delay_signals[0][14]~q ;
wire \fp_functions_0|redist6|delay_signals[0][15]~q ;
wire \fp_functions_0|redist6|delay_signals[0][16]~q ;
wire \fp_functions_0|redist6|delay_signals[0][17]~q ;
wire \fp_functions_0|redist6|delay_signals[0][18]~q ;
wire \fp_functions_0|redist6|delay_signals[0][19]~q ;
wire \fp_functions_0|redist6|delay_signals[0][20]~q ;
wire \fp_functions_0|redist6|delay_signals[0][21]~q ;
wire \fp_functions_0|redist6|delay_signals[0][22]~q ;
wire \fp_functions_0|redist6|delay_signals[0][23]~q ;
wire \fp_functions_0|redist6|delay_signals[0][24]~q ;
wire \fp_functions_0|redist6|delay_signals[0][25]~q ;
wire \fp_functions_0|redist6|delay_signals[0][26]~q ;
wire \fp_functions_0|redist4|delay_signals[0][0]~q ;
wire \fp_functions_0|redist4|delay_signals[0][1]~q ;
wire \fp_functions_0|redist4|delay_signals[0][2]~q ;
wire \fp_functions_0|redist4|delay_signals[0][3]~q ;
wire \fp_functions_0|redist4|delay_signals[0][4]~q ;
wire \fp_functions_0|redist4|delay_signals[0][5]~q ;
wire \fp_functions_0|redist4|delay_signals[0][6]~q ;
wire \fp_functions_0|redist4|delay_signals[0][7]~q ;
wire \fp_functions_0|redist4|delay_signals[0][8]~q ;
wire \fp_functions_0|redist4|delay_signals[0][9]~q ;
wire \fp_functions_0|redist4|delay_signals[0][10]~q ;
wire \fp_functions_0|redist4|delay_signals[0][11]~q ;
wire \fp_functions_0|redist4|delay_signals[0][12]~q ;
wire \fp_functions_0|redist4|delay_signals[0][13]~q ;
wire \fp_functions_0|redist4|delay_signals[0][14]~q ;
wire \fp_functions_0|redist4|delay_signals[0][15]~q ;
wire \fp_functions_0|redist4|delay_signals[0][16]~q ;
wire \fp_functions_0|redist4|delay_signals[0][17]~q ;
wire \fp_functions_0|redist4|delay_signals[0][18]~q ;
wire \fp_functions_0|redist4|delay_signals[0][19]~q ;
wire \fp_functions_0|redist4|delay_signals[0][20]~q ;
wire \fp_functions_0|redist4|delay_signals[0][21]~q ;
wire \fp_functions_0|redist4|delay_signals[0][22]~q ;
wire \fp_functions_0|redist4|delay_signals[0][23]~q ;
wire \fp_functions_0|redist4|delay_signals[0][24]~q ;
wire \fp_functions_0|redist4|delay_signals[0][25]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][0]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][1]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][2]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][3]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][4]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][5]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][6]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][7]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][8]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][9]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][10]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][11]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][12]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][13]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][14]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][15]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][16]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][17]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][18]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][19]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][20]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][21]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][22]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][23]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][24]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][25]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][26]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][0]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][1]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][2]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][3]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][4]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][5]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][6]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][7]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][8]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][9]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][10]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][11]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][12]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][13]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][14]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][15]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][16]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][17]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][18]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][19]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][20]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][21]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][22]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][23]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][24]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][25]~q ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][26]~q ;
wire \fp_functions_0|redist7|delay_signals[0][0]~q ;
wire \fp_functions_0|redist7|delay_signals[0][1]~q ;
wire \fp_functions_0|redist7|delay_signals[0][2]~q ;
wire \fp_functions_0|redist7|delay_signals[0][3]~q ;
wire \fp_functions_0|redist7|delay_signals[0][4]~q ;
wire \fp_functions_0|redist7|delay_signals[0][5]~q ;
wire \fp_functions_0|redist7|delay_signals[0][6]~q ;
wire \fp_functions_0|redist7|delay_signals[0][7]~q ;
wire \fp_functions_0|redist7|delay_signals[0][8]~q ;
wire \fp_functions_0|redist7|delay_signals[0][9]~q ;
wire \fp_functions_0|redist7|delay_signals[0][10]~q ;
wire \fp_functions_0|redist7|delay_signals[0][11]~q ;
wire \fp_functions_0|redist7|delay_signals[0][12]~q ;
wire \fp_functions_0|redist7|delay_signals[0][13]~q ;
wire \fp_functions_0|redist7|delay_signals[0][14]~q ;
wire \fp_functions_0|redist7|delay_signals[0][15]~q ;
wire \fp_functions_0|redist7|delay_signals[0][16]~q ;
wire \fp_functions_0|redist7|delay_signals[0][17]~q ;
wire \fp_functions_0|redist7|delay_signals[0][18]~q ;
wire \fp_functions_0|redist7|delay_signals[0][19]~q ;
wire \fp_functions_0|redist7|delay_signals[0][20]~q ;
wire \fp_functions_0|redist7|delay_signals[0][21]~q ;
wire \fp_functions_0|redist7|delay_signals[0][22]~q ;
wire \fp_functions_0|redist7|delay_signals[0][23]~q ;
wire \fp_functions_0|redist7|delay_signals[0][24]~q ;
wire \fp_functions_0|redist7|delay_signals[0][25]~q ;
wire \fp_functions_0|redist7|delay_signals[0][26]~q ;
wire \fp_functions_0|redist5|delay_signals[0][1]~q ;
wire \fp_functions_0|redist5|delay_signals[0][2]~q ;
wire \fp_functions_0|redist5|delay_signals[0][3]~q ;
wire \fp_functions_0|redist5|delay_signals[0][4]~q ;
wire \fp_functions_0|redist5|delay_signals[0][5]~q ;
wire \fp_functions_0|redist5|delay_signals[0][6]~q ;
wire \fp_functions_0|redist5|delay_signals[0][7]~q ;
wire \fp_functions_0|redist5|delay_signals[0][8]~q ;
wire \fp_functions_0|redist5|delay_signals[0][9]~q ;
wire \fp_functions_0|redist5|delay_signals[0][10]~q ;
wire \fp_functions_0|redist5|delay_signals[0][11]~q ;
wire \fp_functions_0|redist5|delay_signals[0][12]~q ;
wire \fp_functions_0|redist5|delay_signals[0][13]~q ;
wire \fp_functions_0|redist5|delay_signals[0][14]~q ;
wire \fp_functions_0|redist5|delay_signals[0][15]~q ;
wire \fp_functions_0|redist5|delay_signals[0][16]~q ;
wire \fp_functions_0|redist5|delay_signals[0][17]~q ;
wire \fp_functions_0|redist5|delay_signals[0][18]~q ;
wire \fp_functions_0|redist5|delay_signals[0][19]~q ;
wire \fp_functions_0|redist5|delay_signals[0][20]~q ;
wire \fp_functions_0|redist5|delay_signals[0][21]~q ;
wire \fp_functions_0|redist5|delay_signals[0][22]~q ;
wire \fp_functions_0|redist5|delay_signals[0][23]~q ;
wire \fp_functions_0|redist5|delay_signals[0][24]~q ;
wire \fp_functions_0|redist5|delay_signals[0][25]~q ;
wire \fp_functions_0|redist5|delay_signals[0][26]~q ;
wire \fp_functions_0|expSum_uid44_fpMulTest_o[11]~q ;
wire \fp_functions_0|reduce_nor_7~11_combout ;
wire \fp_functions_0|reduce_nor_7~12_combout ;
wire \fp_functions_0|redist11|delay_signals[0][53]~0_combout ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][0]~0_combout ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][0]~0_combout ;
wire \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][0]~0_combout ;
wire \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][0]~0_combout ;

wire [19:0] \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0_PORTBDATAOUT_bus ;
wire [19:0] \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1_PORTBDATAOUT_bus ;
wire [19:0] \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2_PORTBDATAOUT_bus ;
wire [19:0] \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3_PORTBDATAOUT_bus ;
wire [19:0] \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4_PORTBDATAOUT_bus ;
wire [19:0] \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5_PORTBDATAOUT_bus ;
wire [19:0] \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6_PORTBDATAOUT_bus ;
wire [19:0] \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7_PORTBDATAOUT_bus ;
wire [19:0] \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8_PORTBDATAOUT_bus ;
wire [19:0] \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9_PORTBDATAOUT_bus ;
wire [19:0] \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10_PORTBDATAOUT_bus ;
wire [63:0] \fp_functions_0|mult_2~mac_RESULTA_bus ;
wire [63:0] \fp_functions_0|mult_0~mac_RESULTA_bus ;
wire [63:0] \fp_functions_0|mult_1~12_RESULTA_bus ;
wire [63:0] \fp_functions_0|mult_3~mac_RESULTA_bus ;
wire [63:0] \fp_functions_0|mult_3~mac_CHAINOUT_bus ;
wire [19:0] \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11_PORTBDATAOUT_bus ;

assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_wire[0]  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0_PORTBDATAOUT_bus [0];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0~PORTBDATAOUT1  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0_PORTBDATAOUT_bus [1];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0~PORTBDATAOUT2  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0_PORTBDATAOUT_bus [2];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0~PORTBDATAOUT3  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0_PORTBDATAOUT_bus [3];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0~PORTBDATAOUT4  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0_PORTBDATAOUT_bus [4];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0~PORTBDATAOUT5  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0_PORTBDATAOUT_bus [5];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0~PORTBDATAOUT6  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0_PORTBDATAOUT_bus [6];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0~PORTBDATAOUT7  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0_PORTBDATAOUT_bus [7];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0~PORTBDATAOUT8  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0_PORTBDATAOUT_bus [8];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0~PORTBDATAOUT9  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0_PORTBDATAOUT_bus [9];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0~PORTBDATAOUT10  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0_PORTBDATAOUT_bus [10];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0~PORTBDATAOUT11  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0_PORTBDATAOUT_bus [11];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0~PORTBDATAOUT12  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0_PORTBDATAOUT_bus [12];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0~PORTBDATAOUT13  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0_PORTBDATAOUT_bus [13];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0~PORTBDATAOUT14  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0_PORTBDATAOUT_bus [14];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0~PORTBDATAOUT15  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0_PORTBDATAOUT_bus [15];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0~PORTBDATAOUT16  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0_PORTBDATAOUT_bus [16];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0~PORTBDATAOUT17  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0_PORTBDATAOUT_bus [17];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0~PORTBDATAOUT18  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0_PORTBDATAOUT_bus [18];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0~PORTBDATAOUT19  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0_PORTBDATAOUT_bus [19];

assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_wire[1]  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1_PORTBDATAOUT_bus [0];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1~PORTBDATAOUT1  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1_PORTBDATAOUT_bus [1];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1~PORTBDATAOUT2  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1_PORTBDATAOUT_bus [2];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1~PORTBDATAOUT3  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1_PORTBDATAOUT_bus [3];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1~PORTBDATAOUT4  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1_PORTBDATAOUT_bus [4];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1~PORTBDATAOUT5  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1_PORTBDATAOUT_bus [5];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1~PORTBDATAOUT6  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1_PORTBDATAOUT_bus [6];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1~PORTBDATAOUT7  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1_PORTBDATAOUT_bus [7];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1~PORTBDATAOUT8  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1_PORTBDATAOUT_bus [8];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1~PORTBDATAOUT9  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1_PORTBDATAOUT_bus [9];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1~PORTBDATAOUT10  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1_PORTBDATAOUT_bus [10];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1~PORTBDATAOUT11  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1_PORTBDATAOUT_bus [11];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1~PORTBDATAOUT12  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1_PORTBDATAOUT_bus [12];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1~PORTBDATAOUT13  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1_PORTBDATAOUT_bus [13];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1~PORTBDATAOUT14  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1_PORTBDATAOUT_bus [14];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1~PORTBDATAOUT15  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1_PORTBDATAOUT_bus [15];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1~PORTBDATAOUT16  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1_PORTBDATAOUT_bus [16];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1~PORTBDATAOUT17  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1_PORTBDATAOUT_bus [17];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1~PORTBDATAOUT18  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1_PORTBDATAOUT_bus [18];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1~PORTBDATAOUT19  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1_PORTBDATAOUT_bus [19];

assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_wire[2]  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2_PORTBDATAOUT_bus [0];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2~PORTBDATAOUT1  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2_PORTBDATAOUT_bus [1];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2~PORTBDATAOUT2  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2_PORTBDATAOUT_bus [2];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2~PORTBDATAOUT3  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2_PORTBDATAOUT_bus [3];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2~PORTBDATAOUT4  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2_PORTBDATAOUT_bus [4];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2~PORTBDATAOUT5  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2_PORTBDATAOUT_bus [5];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2~PORTBDATAOUT6  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2_PORTBDATAOUT_bus [6];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2~PORTBDATAOUT7  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2_PORTBDATAOUT_bus [7];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2~PORTBDATAOUT8  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2_PORTBDATAOUT_bus [8];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2~PORTBDATAOUT9  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2_PORTBDATAOUT_bus [9];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2~PORTBDATAOUT10  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2_PORTBDATAOUT_bus [10];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2~PORTBDATAOUT11  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2_PORTBDATAOUT_bus [11];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2~PORTBDATAOUT12  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2_PORTBDATAOUT_bus [12];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2~PORTBDATAOUT13  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2_PORTBDATAOUT_bus [13];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2~PORTBDATAOUT14  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2_PORTBDATAOUT_bus [14];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2~PORTBDATAOUT15  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2_PORTBDATAOUT_bus [15];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2~PORTBDATAOUT16  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2_PORTBDATAOUT_bus [16];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2~PORTBDATAOUT17  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2_PORTBDATAOUT_bus [17];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2~PORTBDATAOUT18  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2_PORTBDATAOUT_bus [18];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2~PORTBDATAOUT19  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2_PORTBDATAOUT_bus [19];

assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_wire[3]  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3_PORTBDATAOUT_bus [0];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3~PORTBDATAOUT1  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3_PORTBDATAOUT_bus [1];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3~PORTBDATAOUT2  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3_PORTBDATAOUT_bus [2];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3~PORTBDATAOUT3  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3_PORTBDATAOUT_bus [3];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3~PORTBDATAOUT4  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3_PORTBDATAOUT_bus [4];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3~PORTBDATAOUT5  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3_PORTBDATAOUT_bus [5];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3~PORTBDATAOUT6  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3_PORTBDATAOUT_bus [6];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3~PORTBDATAOUT7  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3_PORTBDATAOUT_bus [7];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3~PORTBDATAOUT8  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3_PORTBDATAOUT_bus [8];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3~PORTBDATAOUT9  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3_PORTBDATAOUT_bus [9];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3~PORTBDATAOUT10  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3_PORTBDATAOUT_bus [10];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3~PORTBDATAOUT11  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3_PORTBDATAOUT_bus [11];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3~PORTBDATAOUT12  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3_PORTBDATAOUT_bus [12];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3~PORTBDATAOUT13  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3_PORTBDATAOUT_bus [13];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3~PORTBDATAOUT14  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3_PORTBDATAOUT_bus [14];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3~PORTBDATAOUT15  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3_PORTBDATAOUT_bus [15];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3~PORTBDATAOUT16  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3_PORTBDATAOUT_bus [16];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3~PORTBDATAOUT17  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3_PORTBDATAOUT_bus [17];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3~PORTBDATAOUT18  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3_PORTBDATAOUT_bus [18];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3~PORTBDATAOUT19  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3_PORTBDATAOUT_bus [19];

assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_wire[4]  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4_PORTBDATAOUT_bus [0];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4~PORTBDATAOUT1  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4_PORTBDATAOUT_bus [1];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4~PORTBDATAOUT2  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4_PORTBDATAOUT_bus [2];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4~PORTBDATAOUT3  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4_PORTBDATAOUT_bus [3];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4~PORTBDATAOUT4  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4_PORTBDATAOUT_bus [4];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4~PORTBDATAOUT5  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4_PORTBDATAOUT_bus [5];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4~PORTBDATAOUT6  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4_PORTBDATAOUT_bus [6];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4~PORTBDATAOUT7  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4_PORTBDATAOUT_bus [7];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4~PORTBDATAOUT8  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4_PORTBDATAOUT_bus [8];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4~PORTBDATAOUT9  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4_PORTBDATAOUT_bus [9];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4~PORTBDATAOUT10  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4_PORTBDATAOUT_bus [10];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4~PORTBDATAOUT11  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4_PORTBDATAOUT_bus [11];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4~PORTBDATAOUT12  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4_PORTBDATAOUT_bus [12];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4~PORTBDATAOUT13  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4_PORTBDATAOUT_bus [13];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4~PORTBDATAOUT14  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4_PORTBDATAOUT_bus [14];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4~PORTBDATAOUT15  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4_PORTBDATAOUT_bus [15];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4~PORTBDATAOUT16  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4_PORTBDATAOUT_bus [16];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4~PORTBDATAOUT17  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4_PORTBDATAOUT_bus [17];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4~PORTBDATAOUT18  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4_PORTBDATAOUT_bus [18];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4~PORTBDATAOUT19  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4_PORTBDATAOUT_bus [19];

assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_wire[5]  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5_PORTBDATAOUT_bus [0];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5~PORTBDATAOUT1  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5_PORTBDATAOUT_bus [1];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5~PORTBDATAOUT2  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5_PORTBDATAOUT_bus [2];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5~PORTBDATAOUT3  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5_PORTBDATAOUT_bus [3];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5~PORTBDATAOUT4  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5_PORTBDATAOUT_bus [4];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5~PORTBDATAOUT5  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5_PORTBDATAOUT_bus [5];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5~PORTBDATAOUT6  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5_PORTBDATAOUT_bus [6];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5~PORTBDATAOUT7  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5_PORTBDATAOUT_bus [7];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5~PORTBDATAOUT8  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5_PORTBDATAOUT_bus [8];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5~PORTBDATAOUT9  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5_PORTBDATAOUT_bus [9];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5~PORTBDATAOUT10  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5_PORTBDATAOUT_bus [10];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5~PORTBDATAOUT11  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5_PORTBDATAOUT_bus [11];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5~PORTBDATAOUT12  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5_PORTBDATAOUT_bus [12];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5~PORTBDATAOUT13  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5_PORTBDATAOUT_bus [13];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5~PORTBDATAOUT14  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5_PORTBDATAOUT_bus [14];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5~PORTBDATAOUT15  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5_PORTBDATAOUT_bus [15];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5~PORTBDATAOUT16  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5_PORTBDATAOUT_bus [16];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5~PORTBDATAOUT17  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5_PORTBDATAOUT_bus [17];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5~PORTBDATAOUT18  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5_PORTBDATAOUT_bus [18];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5~PORTBDATAOUT19  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5_PORTBDATAOUT_bus [19];

assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_wire[6]  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6_PORTBDATAOUT_bus [0];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6~PORTBDATAOUT1  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6_PORTBDATAOUT_bus [1];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6~PORTBDATAOUT2  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6_PORTBDATAOUT_bus [2];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6~PORTBDATAOUT3  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6_PORTBDATAOUT_bus [3];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6~PORTBDATAOUT4  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6_PORTBDATAOUT_bus [4];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6~PORTBDATAOUT5  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6_PORTBDATAOUT_bus [5];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6~PORTBDATAOUT6  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6_PORTBDATAOUT_bus [6];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6~PORTBDATAOUT7  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6_PORTBDATAOUT_bus [7];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6~PORTBDATAOUT8  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6_PORTBDATAOUT_bus [8];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6~PORTBDATAOUT9  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6_PORTBDATAOUT_bus [9];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6~PORTBDATAOUT10  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6_PORTBDATAOUT_bus [10];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6~PORTBDATAOUT11  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6_PORTBDATAOUT_bus [11];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6~PORTBDATAOUT12  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6_PORTBDATAOUT_bus [12];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6~PORTBDATAOUT13  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6_PORTBDATAOUT_bus [13];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6~PORTBDATAOUT14  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6_PORTBDATAOUT_bus [14];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6~PORTBDATAOUT15  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6_PORTBDATAOUT_bus [15];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6~PORTBDATAOUT16  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6_PORTBDATAOUT_bus [16];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6~PORTBDATAOUT17  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6_PORTBDATAOUT_bus [17];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6~PORTBDATAOUT18  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6_PORTBDATAOUT_bus [18];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6~PORTBDATAOUT19  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6_PORTBDATAOUT_bus [19];

assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_wire[7]  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7_PORTBDATAOUT_bus [0];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7~PORTBDATAOUT1  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7_PORTBDATAOUT_bus [1];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7~PORTBDATAOUT2  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7_PORTBDATAOUT_bus [2];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7~PORTBDATAOUT3  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7_PORTBDATAOUT_bus [3];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7~PORTBDATAOUT4  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7_PORTBDATAOUT_bus [4];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7~PORTBDATAOUT5  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7_PORTBDATAOUT_bus [5];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7~PORTBDATAOUT6  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7_PORTBDATAOUT_bus [6];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7~PORTBDATAOUT7  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7_PORTBDATAOUT_bus [7];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7~PORTBDATAOUT8  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7_PORTBDATAOUT_bus [8];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7~PORTBDATAOUT9  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7_PORTBDATAOUT_bus [9];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7~PORTBDATAOUT10  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7_PORTBDATAOUT_bus [10];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7~PORTBDATAOUT11  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7_PORTBDATAOUT_bus [11];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7~PORTBDATAOUT12  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7_PORTBDATAOUT_bus [12];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7~PORTBDATAOUT13  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7_PORTBDATAOUT_bus [13];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7~PORTBDATAOUT14  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7_PORTBDATAOUT_bus [14];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7~PORTBDATAOUT15  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7_PORTBDATAOUT_bus [15];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7~PORTBDATAOUT16  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7_PORTBDATAOUT_bus [16];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7~PORTBDATAOUT17  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7_PORTBDATAOUT_bus [17];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7~PORTBDATAOUT18  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7_PORTBDATAOUT_bus [18];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7~PORTBDATAOUT19  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7_PORTBDATAOUT_bus [19];

assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_wire[8]  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8_PORTBDATAOUT_bus [0];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8~PORTBDATAOUT1  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8_PORTBDATAOUT_bus [1];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8~PORTBDATAOUT2  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8_PORTBDATAOUT_bus [2];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8~PORTBDATAOUT3  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8_PORTBDATAOUT_bus [3];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8~PORTBDATAOUT4  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8_PORTBDATAOUT_bus [4];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8~PORTBDATAOUT5  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8_PORTBDATAOUT_bus [5];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8~PORTBDATAOUT6  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8_PORTBDATAOUT_bus [6];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8~PORTBDATAOUT7  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8_PORTBDATAOUT_bus [7];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8~PORTBDATAOUT8  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8_PORTBDATAOUT_bus [8];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8~PORTBDATAOUT9  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8_PORTBDATAOUT_bus [9];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8~PORTBDATAOUT10  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8_PORTBDATAOUT_bus [10];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8~PORTBDATAOUT11  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8_PORTBDATAOUT_bus [11];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8~PORTBDATAOUT12  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8_PORTBDATAOUT_bus [12];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8~PORTBDATAOUT13  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8_PORTBDATAOUT_bus [13];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8~PORTBDATAOUT14  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8_PORTBDATAOUT_bus [14];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8~PORTBDATAOUT15  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8_PORTBDATAOUT_bus [15];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8~PORTBDATAOUT16  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8_PORTBDATAOUT_bus [16];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8~PORTBDATAOUT17  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8_PORTBDATAOUT_bus [17];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8~PORTBDATAOUT18  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8_PORTBDATAOUT_bus [18];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8~PORTBDATAOUT19  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8_PORTBDATAOUT_bus [19];

assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_wire[9]  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9_PORTBDATAOUT_bus [0];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9~PORTBDATAOUT1  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9_PORTBDATAOUT_bus [1];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9~PORTBDATAOUT2  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9_PORTBDATAOUT_bus [2];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9~PORTBDATAOUT3  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9_PORTBDATAOUT_bus [3];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9~PORTBDATAOUT4  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9_PORTBDATAOUT_bus [4];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9~PORTBDATAOUT5  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9_PORTBDATAOUT_bus [5];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9~PORTBDATAOUT6  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9_PORTBDATAOUT_bus [6];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9~PORTBDATAOUT7  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9_PORTBDATAOUT_bus [7];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9~PORTBDATAOUT8  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9_PORTBDATAOUT_bus [8];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9~PORTBDATAOUT9  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9_PORTBDATAOUT_bus [9];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9~PORTBDATAOUT10  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9_PORTBDATAOUT_bus [10];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9~PORTBDATAOUT11  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9_PORTBDATAOUT_bus [11];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9~PORTBDATAOUT12  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9_PORTBDATAOUT_bus [12];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9~PORTBDATAOUT13  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9_PORTBDATAOUT_bus [13];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9~PORTBDATAOUT14  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9_PORTBDATAOUT_bus [14];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9~PORTBDATAOUT15  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9_PORTBDATAOUT_bus [15];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9~PORTBDATAOUT16  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9_PORTBDATAOUT_bus [16];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9~PORTBDATAOUT17  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9_PORTBDATAOUT_bus [17];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9~PORTBDATAOUT18  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9_PORTBDATAOUT_bus [18];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9~PORTBDATAOUT19  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9_PORTBDATAOUT_bus [19];

assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_wire[10]  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10_PORTBDATAOUT_bus [0];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10~PORTBDATAOUT1  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10_PORTBDATAOUT_bus [1];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10~PORTBDATAOUT2  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10_PORTBDATAOUT_bus [2];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10~PORTBDATAOUT3  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10_PORTBDATAOUT_bus [3];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10~PORTBDATAOUT4  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10_PORTBDATAOUT_bus [4];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10~PORTBDATAOUT5  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10_PORTBDATAOUT_bus [5];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10~PORTBDATAOUT6  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10_PORTBDATAOUT_bus [6];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10~PORTBDATAOUT7  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10_PORTBDATAOUT_bus [7];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10~PORTBDATAOUT8  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10_PORTBDATAOUT_bus [8];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10~PORTBDATAOUT9  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10_PORTBDATAOUT_bus [9];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10~PORTBDATAOUT10  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10_PORTBDATAOUT_bus [10];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10~PORTBDATAOUT11  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10_PORTBDATAOUT_bus [11];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10~PORTBDATAOUT12  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10_PORTBDATAOUT_bus [12];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10~PORTBDATAOUT13  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10_PORTBDATAOUT_bus [13];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10~PORTBDATAOUT14  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10_PORTBDATAOUT_bus [14];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10~PORTBDATAOUT15  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10_PORTBDATAOUT_bus [15];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10~PORTBDATAOUT16  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10_PORTBDATAOUT_bus [16];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10~PORTBDATAOUT17  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10_PORTBDATAOUT_bus [17];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10~PORTBDATAOUT18  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10_PORTBDATAOUT_bus [18];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10~PORTBDATAOUT19  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10_PORTBDATAOUT_bus [19];

assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][0]  = \fp_functions_0|mult_2~mac_RESULTA_bus [0];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][1]  = \fp_functions_0|mult_2~mac_RESULTA_bus [1];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][2]  = \fp_functions_0|mult_2~mac_RESULTA_bus [2];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][3]  = \fp_functions_0|mult_2~mac_RESULTA_bus [3];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][4]  = \fp_functions_0|mult_2~mac_RESULTA_bus [4];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][5]  = \fp_functions_0|mult_2~mac_RESULTA_bus [5];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][6]  = \fp_functions_0|mult_2~mac_RESULTA_bus [6];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][7]  = \fp_functions_0|mult_2~mac_RESULTA_bus [7];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][8]  = \fp_functions_0|mult_2~mac_RESULTA_bus [8];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][9]  = \fp_functions_0|mult_2~mac_RESULTA_bus [9];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][10]  = \fp_functions_0|mult_2~mac_RESULTA_bus [10];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][11]  = \fp_functions_0|mult_2~mac_RESULTA_bus [11];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][12]  = \fp_functions_0|mult_2~mac_RESULTA_bus [12];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][13]  = \fp_functions_0|mult_2~mac_RESULTA_bus [13];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][14]  = \fp_functions_0|mult_2~mac_RESULTA_bus [14];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][15]  = \fp_functions_0|mult_2~mac_RESULTA_bus [15];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][16]  = \fp_functions_0|mult_2~mac_RESULTA_bus [16];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][17]  = \fp_functions_0|mult_2~mac_RESULTA_bus [17];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][18]  = \fp_functions_0|mult_2~mac_RESULTA_bus [18];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][19]  = \fp_functions_0|mult_2~mac_RESULTA_bus [19];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][20]  = \fp_functions_0|mult_2~mac_RESULTA_bus [20];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][21]  = \fp_functions_0|mult_2~mac_RESULTA_bus [21];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][22]  = \fp_functions_0|mult_2~mac_RESULTA_bus [22];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][23]  = \fp_functions_0|mult_2~mac_RESULTA_bus [23];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][24]  = \fp_functions_0|mult_2~mac_RESULTA_bus [24];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][25]  = \fp_functions_0|mult_2~mac_RESULTA_bus [25];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][26]  = \fp_functions_0|mult_2~mac_RESULTA_bus [26];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][27]  = \fp_functions_0|mult_2~mac_RESULTA_bus [27];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][28]  = \fp_functions_0|mult_2~mac_RESULTA_bus [28];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][29]  = \fp_functions_0|mult_2~mac_RESULTA_bus [29];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][30]  = \fp_functions_0|mult_2~mac_RESULTA_bus [30];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][31]  = \fp_functions_0|mult_2~mac_RESULTA_bus [31];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][32]  = \fp_functions_0|mult_2~mac_RESULTA_bus [32];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][33]  = \fp_functions_0|mult_2~mac_RESULTA_bus [33];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][34]  = \fp_functions_0|mult_2~mac_RESULTA_bus [34];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][35]  = \fp_functions_0|mult_2~mac_RESULTA_bus [35];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][36]  = \fp_functions_0|mult_2~mac_RESULTA_bus [36];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][37]  = \fp_functions_0|mult_2~mac_RESULTA_bus [37];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][38]  = \fp_functions_0|mult_2~mac_RESULTA_bus [38];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][39]  = \fp_functions_0|mult_2~mac_RESULTA_bus [39];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][40]  = \fp_functions_0|mult_2~mac_RESULTA_bus [40];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][41]  = \fp_functions_0|mult_2~mac_RESULTA_bus [41];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][42]  = \fp_functions_0|mult_2~mac_RESULTA_bus [42];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][43]  = \fp_functions_0|mult_2~mac_RESULTA_bus [43];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][44]  = \fp_functions_0|mult_2~mac_RESULTA_bus [44];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][45]  = \fp_functions_0|mult_2~mac_RESULTA_bus [45];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][46]  = \fp_functions_0|mult_2~mac_RESULTA_bus [46];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][47]  = \fp_functions_0|mult_2~mac_RESULTA_bus [47];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][48]  = \fp_functions_0|mult_2~mac_RESULTA_bus [48];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][49]  = \fp_functions_0|mult_2~mac_RESULTA_bus [49];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][50]  = \fp_functions_0|mult_2~mac_RESULTA_bus [50];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][51]  = \fp_functions_0|mult_2~mac_RESULTA_bus [51];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][52]  = \fp_functions_0|mult_2~mac_RESULTA_bus [52];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][53]  = \fp_functions_0|mult_2~mac_RESULTA_bus [53];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][54]  = \fp_functions_0|mult_2~mac_RESULTA_bus [54];
assign \fp_functions_0|mult_2~12  = \fp_functions_0|mult_2~mac_RESULTA_bus [55];
assign \fp_functions_0|mult_2~13  = \fp_functions_0|mult_2~mac_RESULTA_bus [56];
assign \fp_functions_0|mult_2~14  = \fp_functions_0|mult_2~mac_RESULTA_bus [57];
assign \fp_functions_0|mult_2~15  = \fp_functions_0|mult_2~mac_RESULTA_bus [58];
assign \fp_functions_0|mult_2~16  = \fp_functions_0|mult_2~mac_RESULTA_bus [59];
assign \fp_functions_0|mult_2~17  = \fp_functions_0|mult_2~mac_RESULTA_bus [60];
assign \fp_functions_0|mult_2~18  = \fp_functions_0|mult_2~mac_RESULTA_bus [61];
assign \fp_functions_0|mult_2~19  = \fp_functions_0|mult_2~mac_RESULTA_bus [62];
assign \fp_functions_0|mult_2~20  = \fp_functions_0|mult_2~mac_RESULTA_bus [63];

assign \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][0]  = \fp_functions_0|mult_0~mac_RESULTA_bus [0];
assign \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][1]  = \fp_functions_0|mult_0~mac_RESULTA_bus [1];
assign \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][2]  = \fp_functions_0|mult_0~mac_RESULTA_bus [2];
assign \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][3]  = \fp_functions_0|mult_0~mac_RESULTA_bus [3];
assign \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][4]  = \fp_functions_0|mult_0~mac_RESULTA_bus [4];
assign \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][5]  = \fp_functions_0|mult_0~mac_RESULTA_bus [5];
assign \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][6]  = \fp_functions_0|mult_0~mac_RESULTA_bus [6];
assign \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][7]  = \fp_functions_0|mult_0~mac_RESULTA_bus [7];
assign \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][8]  = \fp_functions_0|mult_0~mac_RESULTA_bus [8];
assign \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][9]  = \fp_functions_0|mult_0~mac_RESULTA_bus [9];
assign \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][10]  = \fp_functions_0|mult_0~mac_RESULTA_bus [10];
assign \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][11]  = \fp_functions_0|mult_0~mac_RESULTA_bus [11];
assign \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][12]  = \fp_functions_0|mult_0~mac_RESULTA_bus [12];
assign \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][13]  = \fp_functions_0|mult_0~mac_RESULTA_bus [13];
assign \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][14]  = \fp_functions_0|mult_0~mac_RESULTA_bus [14];
assign \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][15]  = \fp_functions_0|mult_0~mac_RESULTA_bus [15];
assign \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][16]  = \fp_functions_0|mult_0~mac_RESULTA_bus [16];
assign \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][17]  = \fp_functions_0|mult_0~mac_RESULTA_bus [17];
assign \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][18]  = \fp_functions_0|mult_0~mac_RESULTA_bus [18];
assign \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][19]  = \fp_functions_0|mult_0~mac_RESULTA_bus [19];
assign \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][20]  = \fp_functions_0|mult_0~mac_RESULTA_bus [20];
assign \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][21]  = \fp_functions_0|mult_0~mac_RESULTA_bus [21];
assign \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][22]  = \fp_functions_0|mult_0~mac_RESULTA_bus [22];
assign \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][23]  = \fp_functions_0|mult_0~mac_RESULTA_bus [23];
assign \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][24]  = \fp_functions_0|mult_0~mac_RESULTA_bus [24];
assign \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][25]  = \fp_functions_0|mult_0~mac_RESULTA_bus [25];
assign \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][26]  = \fp_functions_0|mult_0~mac_RESULTA_bus [26];
assign \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][27]  = \fp_functions_0|mult_0~mac_RESULTA_bus [27];
assign \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][28]  = \fp_functions_0|mult_0~mac_RESULTA_bus [28];
assign \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][29]  = \fp_functions_0|mult_0~mac_RESULTA_bus [29];
assign \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][30]  = \fp_functions_0|mult_0~mac_RESULTA_bus [30];
assign \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][31]  = \fp_functions_0|mult_0~mac_RESULTA_bus [31];
assign \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][32]  = \fp_functions_0|mult_0~mac_RESULTA_bus [32];
assign \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][33]  = \fp_functions_0|mult_0~mac_RESULTA_bus [33];
assign \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][34]  = \fp_functions_0|mult_0~mac_RESULTA_bus [34];
assign \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][35]  = \fp_functions_0|mult_0~mac_RESULTA_bus [35];
assign \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][36]  = \fp_functions_0|mult_0~mac_RESULTA_bus [36];
assign \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][37]  = \fp_functions_0|mult_0~mac_RESULTA_bus [37];
assign \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][38]  = \fp_functions_0|mult_0~mac_RESULTA_bus [38];
assign \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][39]  = \fp_functions_0|mult_0~mac_RESULTA_bus [39];
assign \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][40]  = \fp_functions_0|mult_0~mac_RESULTA_bus [40];
assign \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][41]  = \fp_functions_0|mult_0~mac_RESULTA_bus [41];
assign \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][42]  = \fp_functions_0|mult_0~mac_RESULTA_bus [42];
assign \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][43]  = \fp_functions_0|mult_0~mac_RESULTA_bus [43];
assign \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][44]  = \fp_functions_0|mult_0~mac_RESULTA_bus [44];
assign \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][45]  = \fp_functions_0|mult_0~mac_RESULTA_bus [45];
assign \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][46]  = \fp_functions_0|mult_0~mac_RESULTA_bus [46];
assign \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][47]  = \fp_functions_0|mult_0~mac_RESULTA_bus [47];
assign \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][48]  = \fp_functions_0|mult_0~mac_RESULTA_bus [48];
assign \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][49]  = \fp_functions_0|mult_0~mac_RESULTA_bus [49];
assign \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][50]  = \fp_functions_0|mult_0~mac_RESULTA_bus [50];
assign \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][51]  = \fp_functions_0|mult_0~mac_RESULTA_bus [51];
assign \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][52]  = \fp_functions_0|mult_0~mac_RESULTA_bus [52];
assign \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][53]  = \fp_functions_0|mult_0~mac_RESULTA_bus [53];
assign \fp_functions_0|mult_0~12  = \fp_functions_0|mult_0~mac_RESULTA_bus [54];
assign \fp_functions_0|mult_0~13  = \fp_functions_0|mult_0~mac_RESULTA_bus [55];
assign \fp_functions_0|mult_0~14  = \fp_functions_0|mult_0~mac_RESULTA_bus [56];
assign \fp_functions_0|mult_0~15  = \fp_functions_0|mult_0~mac_RESULTA_bus [57];
assign \fp_functions_0|mult_0~16  = \fp_functions_0|mult_0~mac_RESULTA_bus [58];
assign \fp_functions_0|mult_0~17  = \fp_functions_0|mult_0~mac_RESULTA_bus [59];
assign \fp_functions_0|mult_0~18  = \fp_functions_0|mult_0~mac_RESULTA_bus [60];
assign \fp_functions_0|mult_0~19  = \fp_functions_0|mult_0~mac_RESULTA_bus [61];
assign \fp_functions_0|mult_0~20  = \fp_functions_0|mult_0~mac_RESULTA_bus [62];
assign \fp_functions_0|mult_0~21  = \fp_functions_0|mult_0~mac_RESULTA_bus [63];

assign \fp_functions_0|mult_1~12_resulta  = \fp_functions_0|mult_1~12_RESULTA_bus [0];
assign \fp_functions_0|mult_1~13  = \fp_functions_0|mult_1~12_RESULTA_bus [1];
assign \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][2]  = \fp_functions_0|mult_1~12_RESULTA_bus [2];
assign \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][3]  = \fp_functions_0|mult_1~12_RESULTA_bus [3];
assign \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][4]  = \fp_functions_0|mult_1~12_RESULTA_bus [4];
assign \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][5]  = \fp_functions_0|mult_1~12_RESULTA_bus [5];
assign \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][6]  = \fp_functions_0|mult_1~12_RESULTA_bus [6];
assign \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][7]  = \fp_functions_0|mult_1~12_RESULTA_bus [7];
assign \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][8]  = \fp_functions_0|mult_1~12_RESULTA_bus [8];
assign \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][9]  = \fp_functions_0|mult_1~12_RESULTA_bus [9];
assign \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][10]  = \fp_functions_0|mult_1~12_RESULTA_bus [10];
assign \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][11]  = \fp_functions_0|mult_1~12_RESULTA_bus [11];
assign \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][12]  = \fp_functions_0|mult_1~12_RESULTA_bus [12];
assign \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][13]  = \fp_functions_0|mult_1~12_RESULTA_bus [13];
assign \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][14]  = \fp_functions_0|mult_1~12_RESULTA_bus [14];
assign \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][15]  = \fp_functions_0|mult_1~12_RESULTA_bus [15];
assign \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][16]  = \fp_functions_0|mult_1~12_RESULTA_bus [16];
assign \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][17]  = \fp_functions_0|mult_1~12_RESULTA_bus [17];
assign \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][18]  = \fp_functions_0|mult_1~12_RESULTA_bus [18];
assign \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][19]  = \fp_functions_0|mult_1~12_RESULTA_bus [19];
assign \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][20]  = \fp_functions_0|mult_1~12_RESULTA_bus [20];
assign \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][21]  = \fp_functions_0|mult_1~12_RESULTA_bus [21];
assign \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][22]  = \fp_functions_0|mult_1~12_RESULTA_bus [22];
assign \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][23]  = \fp_functions_0|mult_1~12_RESULTA_bus [23];
assign \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][24]  = \fp_functions_0|mult_1~12_RESULTA_bus [24];
assign \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][25]  = \fp_functions_0|mult_1~12_RESULTA_bus [25];
assign \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][26]  = \fp_functions_0|mult_1~12_RESULTA_bus [26];
assign \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][27]  = \fp_functions_0|mult_1~12_RESULTA_bus [27];
assign \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][28]  = \fp_functions_0|mult_1~12_RESULTA_bus [28];
assign \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][29]  = \fp_functions_0|mult_1~12_RESULTA_bus [29];
assign \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][30]  = \fp_functions_0|mult_1~12_RESULTA_bus [30];
assign \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][31]  = \fp_functions_0|mult_1~12_RESULTA_bus [31];
assign \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][32]  = \fp_functions_0|mult_1~12_RESULTA_bus [32];
assign \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][33]  = \fp_functions_0|mult_1~12_RESULTA_bus [33];
assign \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][34]  = \fp_functions_0|mult_1~12_RESULTA_bus [34];
assign \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][35]  = \fp_functions_0|mult_1~12_RESULTA_bus [35];
assign \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][36]  = \fp_functions_0|mult_1~12_RESULTA_bus [36];
assign \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][37]  = \fp_functions_0|mult_1~12_RESULTA_bus [37];
assign \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][38]  = \fp_functions_0|mult_1~12_RESULTA_bus [38];
assign \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][39]  = \fp_functions_0|mult_1~12_RESULTA_bus [39];
assign \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][40]  = \fp_functions_0|mult_1~12_RESULTA_bus [40];
assign \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][41]  = \fp_functions_0|mult_1~12_RESULTA_bus [41];
assign \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][42]  = \fp_functions_0|mult_1~12_RESULTA_bus [42];
assign \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][43]  = \fp_functions_0|mult_1~12_RESULTA_bus [43];
assign \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][44]  = \fp_functions_0|mult_1~12_RESULTA_bus [44];
assign \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][45]  = \fp_functions_0|mult_1~12_RESULTA_bus [45];
assign \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][46]  = \fp_functions_0|mult_1~12_RESULTA_bus [46];
assign \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][47]  = \fp_functions_0|mult_1~12_RESULTA_bus [47];
assign \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][48]  = \fp_functions_0|mult_1~12_RESULTA_bus [48];
assign \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][49]  = \fp_functions_0|mult_1~12_RESULTA_bus [49];
assign \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][50]  = \fp_functions_0|mult_1~12_RESULTA_bus [50];
assign \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][51]  = \fp_functions_0|mult_1~12_RESULTA_bus [51];
assign \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][52]  = \fp_functions_0|mult_1~12_RESULTA_bus [52];
assign \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][53]  = \fp_functions_0|mult_1~12_RESULTA_bus [53];
assign \fp_functions_0|mult_1~14  = \fp_functions_0|mult_1~12_RESULTA_bus [54];
assign \fp_functions_0|mult_1~15  = \fp_functions_0|mult_1~12_RESULTA_bus [55];
assign \fp_functions_0|mult_1~16  = \fp_functions_0|mult_1~12_RESULTA_bus [56];
assign \fp_functions_0|mult_1~17  = \fp_functions_0|mult_1~12_RESULTA_bus [57];
assign \fp_functions_0|mult_1~18  = \fp_functions_0|mult_1~12_RESULTA_bus [58];
assign \fp_functions_0|mult_1~19  = \fp_functions_0|mult_1~12_RESULTA_bus [59];
assign \fp_functions_0|mult_1~20  = \fp_functions_0|mult_1~12_RESULTA_bus [60];
assign \fp_functions_0|mult_1~21  = \fp_functions_0|mult_1~12_RESULTA_bus [61];
assign \fp_functions_0|mult_1~22  = \fp_functions_0|mult_1~12_RESULTA_bus [62];
assign \fp_functions_0|mult_1~23  = \fp_functions_0|mult_1~12_RESULTA_bus [63];

assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][0]  = \fp_functions_0|mult_3~mac_RESULTA_bus [0];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][1]  = \fp_functions_0|mult_3~mac_RESULTA_bus [1];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][2]  = \fp_functions_0|mult_3~mac_RESULTA_bus [2];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][3]  = \fp_functions_0|mult_3~mac_RESULTA_bus [3];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][4]  = \fp_functions_0|mult_3~mac_RESULTA_bus [4];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][5]  = \fp_functions_0|mult_3~mac_RESULTA_bus [5];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][6]  = \fp_functions_0|mult_3~mac_RESULTA_bus [6];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][7]  = \fp_functions_0|mult_3~mac_RESULTA_bus [7];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][8]  = \fp_functions_0|mult_3~mac_RESULTA_bus [8];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][9]  = \fp_functions_0|mult_3~mac_RESULTA_bus [9];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][10]  = \fp_functions_0|mult_3~mac_RESULTA_bus [10];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][11]  = \fp_functions_0|mult_3~mac_RESULTA_bus [11];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][12]  = \fp_functions_0|mult_3~mac_RESULTA_bus [12];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][13]  = \fp_functions_0|mult_3~mac_RESULTA_bus [13];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][14]  = \fp_functions_0|mult_3~mac_RESULTA_bus [14];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][15]  = \fp_functions_0|mult_3~mac_RESULTA_bus [15];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][16]  = \fp_functions_0|mult_3~mac_RESULTA_bus [16];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][17]  = \fp_functions_0|mult_3~mac_RESULTA_bus [17];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][18]  = \fp_functions_0|mult_3~mac_RESULTA_bus [18];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][19]  = \fp_functions_0|mult_3~mac_RESULTA_bus [19];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][20]  = \fp_functions_0|mult_3~mac_RESULTA_bus [20];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][21]  = \fp_functions_0|mult_3~mac_RESULTA_bus [21];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][22]  = \fp_functions_0|mult_3~mac_RESULTA_bus [22];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][23]  = \fp_functions_0|mult_3~mac_RESULTA_bus [23];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][24]  = \fp_functions_0|mult_3~mac_RESULTA_bus [24];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][25]  = \fp_functions_0|mult_3~mac_RESULTA_bus [25];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][26]  = \fp_functions_0|mult_3~mac_RESULTA_bus [26];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][27]  = \fp_functions_0|mult_3~mac_RESULTA_bus [27];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][28]  = \fp_functions_0|mult_3~mac_RESULTA_bus [28];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][29]  = \fp_functions_0|mult_3~mac_RESULTA_bus [29];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][30]  = \fp_functions_0|mult_3~mac_RESULTA_bus [30];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][31]  = \fp_functions_0|mult_3~mac_RESULTA_bus [31];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][32]  = \fp_functions_0|mult_3~mac_RESULTA_bus [32];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][33]  = \fp_functions_0|mult_3~mac_RESULTA_bus [33];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][34]  = \fp_functions_0|mult_3~mac_RESULTA_bus [34];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][35]  = \fp_functions_0|mult_3~mac_RESULTA_bus [35];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][36]  = \fp_functions_0|mult_3~mac_RESULTA_bus [36];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][37]  = \fp_functions_0|mult_3~mac_RESULTA_bus [37];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][38]  = \fp_functions_0|mult_3~mac_RESULTA_bus [38];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][39]  = \fp_functions_0|mult_3~mac_RESULTA_bus [39];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][40]  = \fp_functions_0|mult_3~mac_RESULTA_bus [40];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][41]  = \fp_functions_0|mult_3~mac_RESULTA_bus [41];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][42]  = \fp_functions_0|mult_3~mac_RESULTA_bus [42];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][43]  = \fp_functions_0|mult_3~mac_RESULTA_bus [43];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][44]  = \fp_functions_0|mult_3~mac_RESULTA_bus [44];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][45]  = \fp_functions_0|mult_3~mac_RESULTA_bus [45];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][46]  = \fp_functions_0|mult_3~mac_RESULTA_bus [46];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][47]  = \fp_functions_0|mult_3~mac_RESULTA_bus [47];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][48]  = \fp_functions_0|mult_3~mac_RESULTA_bus [48];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][49]  = \fp_functions_0|mult_3~mac_RESULTA_bus [49];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][50]  = \fp_functions_0|mult_3~mac_RESULTA_bus [50];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][51]  = \fp_functions_0|mult_3~mac_RESULTA_bus [51];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][52]  = \fp_functions_0|mult_3~mac_RESULTA_bus [52];
assign \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[1][53]  = \fp_functions_0|mult_3~mac_RESULTA_bus [53];
assign \fp_functions_0|mult_3~12  = \fp_functions_0|mult_3~mac_RESULTA_bus [54];
assign \fp_functions_0|mult_3~13  = \fp_functions_0|mult_3~mac_RESULTA_bus [55];
assign \fp_functions_0|mult_3~14  = \fp_functions_0|mult_3~mac_RESULTA_bus [56];
assign \fp_functions_0|mult_3~15  = \fp_functions_0|mult_3~mac_RESULTA_bus [57];
assign \fp_functions_0|mult_3~16  = \fp_functions_0|mult_3~mac_RESULTA_bus [58];
assign \fp_functions_0|mult_3~17  = \fp_functions_0|mult_3~mac_RESULTA_bus [59];
assign \fp_functions_0|mult_3~18  = \fp_functions_0|mult_3~mac_RESULTA_bus [60];
assign \fp_functions_0|mult_3~19  = \fp_functions_0|mult_3~mac_RESULTA_bus [61];
assign \fp_functions_0|mult_3~20  = \fp_functions_0|mult_3~mac_RESULTA_bus [62];
assign \fp_functions_0|mult_3~21  = \fp_functions_0|mult_3~mac_RESULTA_bus [63];

assign \fp_functions_0|mult_3~86  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [0];
assign \fp_functions_0|mult_3~87  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [1];
assign \fp_functions_0|mult_3~88  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [2];
assign \fp_functions_0|mult_3~89  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [3];
assign \fp_functions_0|mult_3~90  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [4];
assign \fp_functions_0|mult_3~91  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [5];
assign \fp_functions_0|mult_3~92  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [6];
assign \fp_functions_0|mult_3~93  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [7];
assign \fp_functions_0|mult_3~94  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [8];
assign \fp_functions_0|mult_3~95  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [9];
assign \fp_functions_0|mult_3~96  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [10];
assign \fp_functions_0|mult_3~97  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [11];
assign \fp_functions_0|mult_3~98  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [12];
assign \fp_functions_0|mult_3~99  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [13];
assign \fp_functions_0|mult_3~100  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [14];
assign \fp_functions_0|mult_3~101  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [15];
assign \fp_functions_0|mult_3~102  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [16];
assign \fp_functions_0|mult_3~103  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [17];
assign \fp_functions_0|mult_3~104  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [18];
assign \fp_functions_0|mult_3~105  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [19];
assign \fp_functions_0|mult_3~106  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [20];
assign \fp_functions_0|mult_3~107  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [21];
assign \fp_functions_0|mult_3~108  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [22];
assign \fp_functions_0|mult_3~109  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [23];
assign \fp_functions_0|mult_3~110  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [24];
assign \fp_functions_0|mult_3~111  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [25];
assign \fp_functions_0|mult_3~112  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [26];
assign \fp_functions_0|mult_3~113  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [27];
assign \fp_functions_0|mult_3~114  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [28];
assign \fp_functions_0|mult_3~115  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [29];
assign \fp_functions_0|mult_3~116  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [30];
assign \fp_functions_0|mult_3~117  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [31];
assign \fp_functions_0|mult_3~118  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [32];
assign \fp_functions_0|mult_3~119  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [33];
assign \fp_functions_0|mult_3~120  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [34];
assign \fp_functions_0|mult_3~121  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [35];
assign \fp_functions_0|mult_3~122  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [36];
assign \fp_functions_0|mult_3~123  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [37];
assign \fp_functions_0|mult_3~124  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [38];
assign \fp_functions_0|mult_3~125  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [39];
assign \fp_functions_0|mult_3~126  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [40];
assign \fp_functions_0|mult_3~127  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [41];
assign \fp_functions_0|mult_3~128  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [42];
assign \fp_functions_0|mult_3~129  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [43];
assign \fp_functions_0|mult_3~130  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [44];
assign \fp_functions_0|mult_3~131  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [45];
assign \fp_functions_0|mult_3~132  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [46];
assign \fp_functions_0|mult_3~133  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [47];
assign \fp_functions_0|mult_3~134  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [48];
assign \fp_functions_0|mult_3~135  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [49];
assign \fp_functions_0|mult_3~136  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [50];
assign \fp_functions_0|mult_3~137  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [51];
assign \fp_functions_0|mult_3~138  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [52];
assign \fp_functions_0|mult_3~139  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [53];
assign \fp_functions_0|mult_3~140  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [54];
assign \fp_functions_0|mult_3~141  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [55];
assign \fp_functions_0|mult_3~142  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [56];
assign \fp_functions_0|mult_3~143  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [57];
assign \fp_functions_0|mult_3~144  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [58];
assign \fp_functions_0|mult_3~145  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [59];
assign \fp_functions_0|mult_3~146  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [60];
assign \fp_functions_0|mult_3~147  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [61];
assign \fp_functions_0|mult_3~148  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [62];
assign \fp_functions_0|mult_3~149  = \fp_functions_0|mult_3~mac_CHAINOUT_bus [63];

assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_wire[11]  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11_PORTBDATAOUT_bus [0];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11~PORTBDATAOUT1  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11_PORTBDATAOUT_bus [1];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11~PORTBDATAOUT2  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11_PORTBDATAOUT_bus [2];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11~PORTBDATAOUT3  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11_PORTBDATAOUT_bus [3];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11~PORTBDATAOUT4  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11_PORTBDATAOUT_bus [4];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11~PORTBDATAOUT5  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11_PORTBDATAOUT_bus [5];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11~PORTBDATAOUT6  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11_PORTBDATAOUT_bus [6];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11~PORTBDATAOUT7  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11_PORTBDATAOUT_bus [7];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11~PORTBDATAOUT8  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11_PORTBDATAOUT_bus [8];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11~PORTBDATAOUT9  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11_PORTBDATAOUT_bus [9];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11~PORTBDATAOUT10  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11_PORTBDATAOUT_bus [10];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11~PORTBDATAOUT11  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11_PORTBDATAOUT_bus [11];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11~PORTBDATAOUT12  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11_PORTBDATAOUT_bus [12];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11~PORTBDATAOUT13  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11_PORTBDATAOUT_bus [13];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11~PORTBDATAOUT14  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11_PORTBDATAOUT_bus [14];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11~PORTBDATAOUT15  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11_PORTBDATAOUT_bus [15];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11~PORTBDATAOUT16  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11_PORTBDATAOUT_bus [16];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11~PORTBDATAOUT17  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11_PORTBDATAOUT_bus [17];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11~PORTBDATAOUT18  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11_PORTBDATAOUT_bus [18];
assign \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11~PORTBDATAOUT19  = \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11_PORTBDATAOUT_bus [19];

twentynm_lcell_comb \fp_functions_0|add_7~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist9|delay_signals[0][14]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_7~6_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_7~1_sumout ),
	.cout(),
	.shareout());
defparam \fp_functions_0|add_7~1 .extended_lut = "off";
defparam \fp_functions_0|add_7~1 .lut_mask = 64'h00000000000000FF;
defparam \fp_functions_0|add_7~1 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_8~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist9|delay_signals[0][14]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_8~6_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_8~1_sumout ),
	.cout(),
	.shareout());
defparam \fp_functions_0|add_8~1 .extended_lut = "off";
defparam \fp_functions_0|add_8~1 .lut_mask = 64'h0000FFFF0000FF00;
defparam \fp_functions_0|add_8~1 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~254_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~1_sumout ),
	.cout(\fp_functions_0|add_6~2 ),
	.shareout());
defparam \fp_functions_0|add_6~1 .extended_lut = "off";
defparam \fp_functions_0|add_6~1 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~1 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_7~6 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist9|delay_signals[0][14]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_7~10_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fp_functions_0|add_7~6_cout ),
	.shareout());
defparam \fp_functions_0|add_7~6 .extended_lut = "off";
defparam \fp_functions_0|add_7~6 .lut_mask = 64'h00000000000000FF;
defparam \fp_functions_0|add_7~6 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_8~6 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist9|delay_signals[0][14]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_8~10_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fp_functions_0|add_8~6_cout ),
	.shareout());
defparam \fp_functions_0|add_8~6 .extended_lut = "off";
defparam \fp_functions_0|add_8~6 .lut_mask = 64'h0000FFFF0000FF00;
defparam \fp_functions_0|add_8~6 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~5_sumout ),
	.cout(\fp_functions_0|add_6~6 ),
	.shareout());
defparam \fp_functions_0|add_6~5 .extended_lut = "off";
defparam \fp_functions_0|add_6~5 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~5 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~9_sumout ),
	.cout(\fp_functions_0|add_6~10 ),
	.shareout());
defparam \fp_functions_0|add_6~9 .extended_lut = "off";
defparam \fp_functions_0|add_6~9 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~9 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~13_sumout ),
	.cout(\fp_functions_0|add_6~14 ),
	.shareout());
defparam \fp_functions_0|add_6~13 .extended_lut = "off";
defparam \fp_functions_0|add_6~13 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~13 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~17_sumout ),
	.cout(\fp_functions_0|add_6~18 ),
	.shareout());
defparam \fp_functions_0|add_6~17 .extended_lut = "off";
defparam \fp_functions_0|add_6~17 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~17 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~21_sumout ),
	.cout(\fp_functions_0|add_6~22 ),
	.shareout());
defparam \fp_functions_0|add_6~21 .extended_lut = "off";
defparam \fp_functions_0|add_6~21 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~21 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~25_sumout ),
	.cout(\fp_functions_0|add_6~26 ),
	.shareout());
defparam \fp_functions_0|add_6~25 .extended_lut = "off";
defparam \fp_functions_0|add_6~25 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~25 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~29_sumout ),
	.cout(\fp_functions_0|add_6~30 ),
	.shareout());
defparam \fp_functions_0|add_6~29 .extended_lut = "off";
defparam \fp_functions_0|add_6~29 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~29 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~33_sumout ),
	.cout(\fp_functions_0|add_6~34 ),
	.shareout());
defparam \fp_functions_0|add_6~33 .extended_lut = "off";
defparam \fp_functions_0|add_6~33 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~33 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~37_sumout ),
	.cout(\fp_functions_0|add_6~38 ),
	.shareout());
defparam \fp_functions_0|add_6~37 .extended_lut = "off";
defparam \fp_functions_0|add_6~37 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~37 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][11]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~41_sumout ),
	.cout(\fp_functions_0|add_6~42 ),
	.shareout());
defparam \fp_functions_0|add_6~41 .extended_lut = "off";
defparam \fp_functions_0|add_6~41 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~41 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~45_sumout ),
	.cout(\fp_functions_0|add_6~46 ),
	.shareout());
defparam \fp_functions_0|add_6~45 .extended_lut = "off";
defparam \fp_functions_0|add_6~45 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~45 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][13]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~49_sumout ),
	.cout(\fp_functions_0|add_6~50 ),
	.shareout());
defparam \fp_functions_0|add_6~49 .extended_lut = "off";
defparam \fp_functions_0|add_6~49 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~49 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][14]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~53_sumout ),
	.cout(\fp_functions_0|add_6~54 ),
	.shareout());
defparam \fp_functions_0|add_6~53 .extended_lut = "off";
defparam \fp_functions_0|add_6~53 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~53 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][15]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~57_sumout ),
	.cout(\fp_functions_0|add_6~58 ),
	.shareout());
defparam \fp_functions_0|add_6~57 .extended_lut = "off";
defparam \fp_functions_0|add_6~57 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~57 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][16]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~61_sumout ),
	.cout(\fp_functions_0|add_6~62 ),
	.shareout());
defparam \fp_functions_0|add_6~61 .extended_lut = "off";
defparam \fp_functions_0|add_6~61 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~61 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][17]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~65_sumout ),
	.cout(\fp_functions_0|add_6~66 ),
	.shareout());
defparam \fp_functions_0|add_6~65 .extended_lut = "off";
defparam \fp_functions_0|add_6~65 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~65 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][18]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~69_sumout ),
	.cout(\fp_functions_0|add_6~70 ),
	.shareout());
defparam \fp_functions_0|add_6~69 .extended_lut = "off";
defparam \fp_functions_0|add_6~69 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~69 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~73 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][19]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~73_sumout ),
	.cout(\fp_functions_0|add_6~74 ),
	.shareout());
defparam \fp_functions_0|add_6~73 .extended_lut = "off";
defparam \fp_functions_0|add_6~73 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~73 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~77 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][20]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~74 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~77_sumout ),
	.cout(\fp_functions_0|add_6~78 ),
	.shareout());
defparam \fp_functions_0|add_6~77 .extended_lut = "off";
defparam \fp_functions_0|add_6~77 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~77 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~81 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][21]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~78 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~81_sumout ),
	.cout(\fp_functions_0|add_6~82 ),
	.shareout());
defparam \fp_functions_0|add_6~81 .extended_lut = "off";
defparam \fp_functions_0|add_6~81 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~81 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~85 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][22]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~82 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~85_sumout ),
	.cout(\fp_functions_0|add_6~86 ),
	.shareout());
defparam \fp_functions_0|add_6~85 .extended_lut = "off";
defparam \fp_functions_0|add_6~85 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~85 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~89 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][23]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~86 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~89_sumout ),
	.cout(\fp_functions_0|add_6~90 ),
	.shareout());
defparam \fp_functions_0|add_6~89 .extended_lut = "off";
defparam \fp_functions_0|add_6~89 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~89 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~93 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][24]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~90 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~93_sumout ),
	.cout(\fp_functions_0|add_6~94 ),
	.shareout());
defparam \fp_functions_0|add_6~93 .extended_lut = "off";
defparam \fp_functions_0|add_6~93 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~93 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~97 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][25]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~94 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~97_sumout ),
	.cout(\fp_functions_0|add_6~98 ),
	.shareout());
defparam \fp_functions_0|add_6~97 .extended_lut = "off";
defparam \fp_functions_0|add_6~97 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~97 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~101 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][26]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~98 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~101_sumout ),
	.cout(\fp_functions_0|add_6~102 ),
	.shareout());
defparam \fp_functions_0|add_6~101 .extended_lut = "off";
defparam \fp_functions_0|add_6~101 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~101 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~105 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][27]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~102 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~105_sumout ),
	.cout(\fp_functions_0|add_6~106 ),
	.shareout());
defparam \fp_functions_0|add_6~105 .extended_lut = "off";
defparam \fp_functions_0|add_6~105 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~105 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~109 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][28]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~106 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~109_sumout ),
	.cout(\fp_functions_0|add_6~110 ),
	.shareout());
defparam \fp_functions_0|add_6~109 .extended_lut = "off";
defparam \fp_functions_0|add_6~109 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~109 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~113 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][29]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~110 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~113_sumout ),
	.cout(\fp_functions_0|add_6~114 ),
	.shareout());
defparam \fp_functions_0|add_6~113 .extended_lut = "off";
defparam \fp_functions_0|add_6~113 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~113 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~117 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][30]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~114 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~117_sumout ),
	.cout(\fp_functions_0|add_6~118 ),
	.shareout());
defparam \fp_functions_0|add_6~117 .extended_lut = "off";
defparam \fp_functions_0|add_6~117 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~117 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~121 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][31]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~118 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~121_sumout ),
	.cout(\fp_functions_0|add_6~122 ),
	.shareout());
defparam \fp_functions_0|add_6~121 .extended_lut = "off";
defparam \fp_functions_0|add_6~121 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~121 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~125 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][32]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~122 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~125_sumout ),
	.cout(\fp_functions_0|add_6~126 ),
	.shareout());
defparam \fp_functions_0|add_6~125 .extended_lut = "off";
defparam \fp_functions_0|add_6~125 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~125 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~129 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][33]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~126 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~129_sumout ),
	.cout(\fp_functions_0|add_6~130 ),
	.shareout());
defparam \fp_functions_0|add_6~129 .extended_lut = "off";
defparam \fp_functions_0|add_6~129 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~129 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~133 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][34]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~130 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~133_sumout ),
	.cout(\fp_functions_0|add_6~134 ),
	.shareout());
defparam \fp_functions_0|add_6~133 .extended_lut = "off";
defparam \fp_functions_0|add_6~133 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~133 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~137 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][35]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~134 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~137_sumout ),
	.cout(\fp_functions_0|add_6~138 ),
	.shareout());
defparam \fp_functions_0|add_6~137 .extended_lut = "off";
defparam \fp_functions_0|add_6~137 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~137 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~141 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][36]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~138 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~141_sumout ),
	.cout(\fp_functions_0|add_6~142 ),
	.shareout());
defparam \fp_functions_0|add_6~141 .extended_lut = "off";
defparam \fp_functions_0|add_6~141 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~141 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~145 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][37]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~142 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~145_sumout ),
	.cout(\fp_functions_0|add_6~146 ),
	.shareout());
defparam \fp_functions_0|add_6~145 .extended_lut = "off";
defparam \fp_functions_0|add_6~145 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~145 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~149 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][38]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~146 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~149_sumout ),
	.cout(\fp_functions_0|add_6~150 ),
	.shareout());
defparam \fp_functions_0|add_6~149 .extended_lut = "off";
defparam \fp_functions_0|add_6~149 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~149 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~153 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][39]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~150 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~153_sumout ),
	.cout(\fp_functions_0|add_6~154 ),
	.shareout());
defparam \fp_functions_0|add_6~153 .extended_lut = "off";
defparam \fp_functions_0|add_6~153 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~153 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~157 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][40]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~154 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~157_sumout ),
	.cout(\fp_functions_0|add_6~158 ),
	.shareout());
defparam \fp_functions_0|add_6~157 .extended_lut = "off";
defparam \fp_functions_0|add_6~157 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~157 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~161 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][41]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~158 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~161_sumout ),
	.cout(\fp_functions_0|add_6~162 ),
	.shareout());
defparam \fp_functions_0|add_6~161 .extended_lut = "off";
defparam \fp_functions_0|add_6~161 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~161 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~165 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][42]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~162 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~165_sumout ),
	.cout(\fp_functions_0|add_6~166 ),
	.shareout());
defparam \fp_functions_0|add_6~165 .extended_lut = "off";
defparam \fp_functions_0|add_6~165 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~165 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~169 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][43]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~166 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~169_sumout ),
	.cout(\fp_functions_0|add_6~170 ),
	.shareout());
defparam \fp_functions_0|add_6~169 .extended_lut = "off";
defparam \fp_functions_0|add_6~169 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~169 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~173 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][44]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~170 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~173_sumout ),
	.cout(\fp_functions_0|add_6~174 ),
	.shareout());
defparam \fp_functions_0|add_6~173 .extended_lut = "off";
defparam \fp_functions_0|add_6~173 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~173 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~177 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][45]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~174 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~177_sumout ),
	.cout(\fp_functions_0|add_6~178 ),
	.shareout());
defparam \fp_functions_0|add_6~177 .extended_lut = "off";
defparam \fp_functions_0|add_6~177 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~177 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~181 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][46]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~178 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~181_sumout ),
	.cout(\fp_functions_0|add_6~182 ),
	.shareout());
defparam \fp_functions_0|add_6~181 .extended_lut = "off";
defparam \fp_functions_0|add_6~181 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~181 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~185 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][47]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~182 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~185_sumout ),
	.cout(\fp_functions_0|add_6~186 ),
	.shareout());
defparam \fp_functions_0|add_6~185 .extended_lut = "off";
defparam \fp_functions_0|add_6~185 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~185 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~189 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][48]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~186 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~189_sumout ),
	.cout(\fp_functions_0|add_6~190 ),
	.shareout());
defparam \fp_functions_0|add_6~189 .extended_lut = "off";
defparam \fp_functions_0|add_6~189 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~189 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~193 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][49]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~190 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~193_sumout ),
	.cout(\fp_functions_0|add_6~194 ),
	.shareout());
defparam \fp_functions_0|add_6~193 .extended_lut = "off";
defparam \fp_functions_0|add_6~193 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~193 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~197 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][50]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~194 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~197_sumout ),
	.cout(\fp_functions_0|add_6~198 ),
	.shareout());
defparam \fp_functions_0|add_6~197 .extended_lut = "off";
defparam \fp_functions_0|add_6~197 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~197 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~201 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][51]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~198 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~201_sumout ),
	.cout(\fp_functions_0|add_6~202 ),
	.shareout());
defparam \fp_functions_0|add_6~201 .extended_lut = "off";
defparam \fp_functions_0|add_6~201 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~201 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~205 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][52]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~202 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~205_sumout ),
	.cout(\fp_functions_0|add_6~206 ),
	.shareout());
defparam \fp_functions_0|add_6~205 .extended_lut = "off";
defparam \fp_functions_0|add_6~205 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~205 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~209 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][53]~q ),
	.datae(gnd),
	.dataf(!\fp_functions_0|redist13|delay_signals[0][0]~q ),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~206 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~209_sumout ),
	.cout(\fp_functions_0|add_6~210 ),
	.shareout());
defparam \fp_functions_0|add_6~209 .extended_lut = "off";
defparam \fp_functions_0|add_6~209 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_6~209 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~213 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][54]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~210 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~213_sumout ),
	.cout(\fp_functions_0|add_6~214 ),
	.shareout());
defparam \fp_functions_0|add_6~213 .extended_lut = "off";
defparam \fp_functions_0|add_6~213 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~213 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~217 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][55]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~214 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~217_sumout ),
	.cout(\fp_functions_0|add_6~218 ),
	.shareout());
defparam \fp_functions_0|add_6~217 .extended_lut = "off";
defparam \fp_functions_0|add_6~217 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~217 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~221 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][56]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~218 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~221_sumout ),
	.cout(\fp_functions_0|add_6~222 ),
	.shareout());
defparam \fp_functions_0|add_6~221 .extended_lut = "off";
defparam \fp_functions_0|add_6~221 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~221 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~225 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][57]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~222 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~225_sumout ),
	.cout(\fp_functions_0|add_6~226 ),
	.shareout());
defparam \fp_functions_0|add_6~225 .extended_lut = "off";
defparam \fp_functions_0|add_6~225 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~225 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~229 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][58]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~226 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~229_sumout ),
	.cout(\fp_functions_0|add_6~230 ),
	.shareout());
defparam \fp_functions_0|add_6~229 .extended_lut = "off";
defparam \fp_functions_0|add_6~229 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~229 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~233 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][59]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~230 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~233_sumout ),
	.cout(\fp_functions_0|add_6~234 ),
	.shareout());
defparam \fp_functions_0|add_6~233 .extended_lut = "off";
defparam \fp_functions_0|add_6~233 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~233 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~237 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][60]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~234 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~237_sumout ),
	.cout(\fp_functions_0|add_6~238 ),
	.shareout());
defparam \fp_functions_0|add_6~237 .extended_lut = "off";
defparam \fp_functions_0|add_6~237 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~237 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~241 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][61]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~238 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~241_sumout ),
	.cout(\fp_functions_0|add_6~242 ),
	.shareout());
defparam \fp_functions_0|add_6~241 .extended_lut = "off";
defparam \fp_functions_0|add_6~241 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~241 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~245 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][62]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~242 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~245_sumout ),
	.cout(\fp_functions_0|add_6~246 ),
	.shareout());
defparam \fp_functions_0|add_6~245 .extended_lut = "off";
defparam \fp_functions_0|add_6~245 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~245 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~249 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][63]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~246 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~249_sumout ),
	.cout(\fp_functions_0|add_6~250 ),
	.shareout());
defparam \fp_functions_0|add_6~249 .extended_lut = "off";
defparam \fp_functions_0|add_6~249 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~249 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~254 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][0]~q ),
	.datae(gnd),
	.dataf(!\fp_functions_0|roundBit_uid65_fpMulTest_delay|delay_signals[0][0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fp_functions_0|add_6~254_cout ),
	.shareout());
defparam \fp_functions_0|add_6~254 .extended_lut = "off";
defparam \fp_functions_0|add_6~254 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_6~254 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~257 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][66]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~262 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~257_sumout ),
	.cout(),
	.shareout());
defparam \fp_functions_0|add_6~257 .extended_lut = "off";
defparam \fp_functions_0|add_6~257 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~257 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_7~10 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist9|delay_signals[0][13]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_7~14_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fp_functions_0|add_7~10_cout ),
	.shareout());
defparam \fp_functions_0|add_7~10 .extended_lut = "off";
defparam \fp_functions_0|add_7~10 .lut_mask = 64'h00000000000000FF;
defparam \fp_functions_0|add_7~10 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_8~10 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist9|delay_signals[0][13]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_8~14_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fp_functions_0|add_8~10_cout ),
	.shareout());
defparam \fp_functions_0|add_8~10 .extended_lut = "off";
defparam \fp_functions_0|add_8~10 .lut_mask = 64'h0000FFFF0000FF00;
defparam \fp_functions_0|add_8~10 .shared_arith = "off";

dffeas \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[1] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][52]~q ),
	.asdata(\fp_functions_0|redist1|delay_signals[0][53]~q ),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\fp_functions_0|redist1|delay_signals[0][105]~q ),
	.ena(en[0]),
	.q(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[1]~q ),
	.prn(vcc));
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[1] .is_wysiwyg = "true";
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[1] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|add_6~261 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][66]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~266 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~261_sumout ),
	.cout(\fp_functions_0|add_6~262 ),
	.shareout());
defparam \fp_functions_0|add_6~261 .extended_lut = "off";
defparam \fp_functions_0|add_6~261 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~261 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_7~14 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist9|delay_signals[0][12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_7~18_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fp_functions_0|add_7~14_cout ),
	.shareout());
defparam \fp_functions_0|add_7~14 .extended_lut = "off";
defparam \fp_functions_0|add_7~14 .lut_mask = 64'h00000000000000FF;
defparam \fp_functions_0|add_7~14 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_8~14 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist9|delay_signals[0][12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_8~18_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fp_functions_0|add_8~14_cout ),
	.shareout());
defparam \fp_functions_0|add_8~14 .extended_lut = "off";
defparam \fp_functions_0|add_8~14 .lut_mask = 64'h0000FFFF0000FF00;
defparam \fp_functions_0|add_8~14 .shared_arith = "off";

dffeas \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[2] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][53]~q ),
	.asdata(\fp_functions_0|redist1|delay_signals[0][54]~q ),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\fp_functions_0|redist1|delay_signals[0][105]~q ),
	.ena(en[0]),
	.q(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[2]~q ),
	.prn(vcc));
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[2] .is_wysiwyg = "true";
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[2] .power_up = "low";

dffeas \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[3] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][54]~q ),
	.asdata(\fp_functions_0|redist1|delay_signals[0][55]~q ),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\fp_functions_0|redist1|delay_signals[0][105]~q ),
	.ena(en[0]),
	.q(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[3]~q ),
	.prn(vcc));
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[3] .is_wysiwyg = "true";
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[3] .power_up = "low";

dffeas \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[4] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][55]~q ),
	.asdata(\fp_functions_0|redist1|delay_signals[0][56]~q ),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\fp_functions_0|redist1|delay_signals[0][105]~q ),
	.ena(en[0]),
	.q(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[4]~q ),
	.prn(vcc));
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[4] .is_wysiwyg = "true";
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[4] .power_up = "low";

dffeas \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[5] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][56]~q ),
	.asdata(\fp_functions_0|redist1|delay_signals[0][57]~q ),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\fp_functions_0|redist1|delay_signals[0][105]~q ),
	.ena(en[0]),
	.q(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[5]~q ),
	.prn(vcc));
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[5] .is_wysiwyg = "true";
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[5] .power_up = "low";

dffeas \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[6] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][57]~q ),
	.asdata(\fp_functions_0|redist1|delay_signals[0][58]~q ),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\fp_functions_0|redist1|delay_signals[0][105]~q ),
	.ena(en[0]),
	.q(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[6]~q ),
	.prn(vcc));
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[6] .is_wysiwyg = "true";
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[6] .power_up = "low";

dffeas \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[7] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][58]~q ),
	.asdata(\fp_functions_0|redist1|delay_signals[0][59]~q ),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\fp_functions_0|redist1|delay_signals[0][105]~q ),
	.ena(en[0]),
	.q(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[7]~q ),
	.prn(vcc));
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[7] .is_wysiwyg = "true";
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[7] .power_up = "low";

dffeas \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[8] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][59]~q ),
	.asdata(\fp_functions_0|redist1|delay_signals[0][60]~q ),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\fp_functions_0|redist1|delay_signals[0][105]~q ),
	.ena(en[0]),
	.q(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[8]~q ),
	.prn(vcc));
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[8] .is_wysiwyg = "true";
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[8] .power_up = "low";

dffeas \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[9] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][60]~q ),
	.asdata(\fp_functions_0|redist1|delay_signals[0][61]~q ),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\fp_functions_0|redist1|delay_signals[0][105]~q ),
	.ena(en[0]),
	.q(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[9]~q ),
	.prn(vcc));
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[9] .is_wysiwyg = "true";
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[9] .power_up = "low";

dffeas \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[10] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][61]~q ),
	.asdata(\fp_functions_0|redist1|delay_signals[0][62]~q ),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\fp_functions_0|redist1|delay_signals[0][105]~q ),
	.ena(en[0]),
	.q(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[10]~q ),
	.prn(vcc));
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[10] .is_wysiwyg = "true";
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[10] .power_up = "low";

dffeas \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[11] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][62]~q ),
	.asdata(\fp_functions_0|redist1|delay_signals[0][63]~q ),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\fp_functions_0|redist1|delay_signals[0][105]~q ),
	.ena(en[0]),
	.q(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[11]~q ),
	.prn(vcc));
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[11] .is_wysiwyg = "true";
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[11] .power_up = "low";

dffeas \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[12] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][63]~q ),
	.asdata(\fp_functions_0|redist1|delay_signals[0][64]~q ),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\fp_functions_0|redist1|delay_signals[0][105]~q ),
	.ena(en[0]),
	.q(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[12]~q ),
	.prn(vcc));
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[12] .is_wysiwyg = "true";
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[12] .power_up = "low";

dffeas \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[13] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][64]~q ),
	.asdata(\fp_functions_0|redist1|delay_signals[0][65]~q ),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\fp_functions_0|redist1|delay_signals[0][105]~q ),
	.ena(en[0]),
	.q(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[13]~q ),
	.prn(vcc));
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[13] .is_wysiwyg = "true";
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[13] .power_up = "low";

dffeas \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[14] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][65]~q ),
	.asdata(\fp_functions_0|redist1|delay_signals[0][66]~q ),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\fp_functions_0|redist1|delay_signals[0][105]~q ),
	.ena(en[0]),
	.q(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[14]~q ),
	.prn(vcc));
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[14] .is_wysiwyg = "true";
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[14] .power_up = "low";

dffeas \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[15] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][66]~q ),
	.asdata(\fp_functions_0|redist1|delay_signals[0][67]~q ),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\fp_functions_0|redist1|delay_signals[0][105]~q ),
	.ena(en[0]),
	.q(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[15]~q ),
	.prn(vcc));
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[15] .is_wysiwyg = "true";
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[15] .power_up = "low";

dffeas \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[16] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][67]~q ),
	.asdata(\fp_functions_0|redist1|delay_signals[0][68]~q ),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\fp_functions_0|redist1|delay_signals[0][105]~q ),
	.ena(en[0]),
	.q(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[16]~q ),
	.prn(vcc));
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[16] .is_wysiwyg = "true";
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[16] .power_up = "low";

dffeas \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[17] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][68]~q ),
	.asdata(\fp_functions_0|redist1|delay_signals[0][69]~q ),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\fp_functions_0|redist1|delay_signals[0][105]~q ),
	.ena(en[0]),
	.q(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[17]~q ),
	.prn(vcc));
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[17] .is_wysiwyg = "true";
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[17] .power_up = "low";

dffeas \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[18] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][69]~q ),
	.asdata(\fp_functions_0|redist1|delay_signals[0][70]~q ),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\fp_functions_0|redist1|delay_signals[0][105]~q ),
	.ena(en[0]),
	.q(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[18]~q ),
	.prn(vcc));
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[18] .is_wysiwyg = "true";
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[18] .power_up = "low";

dffeas \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[19] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][70]~q ),
	.asdata(\fp_functions_0|redist1|delay_signals[0][71]~q ),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\fp_functions_0|redist1|delay_signals[0][105]~q ),
	.ena(en[0]),
	.q(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[19]~q ),
	.prn(vcc));
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[19] .is_wysiwyg = "true";
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[19] .power_up = "low";

dffeas \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[20] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][71]~q ),
	.asdata(\fp_functions_0|redist1|delay_signals[0][72]~q ),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\fp_functions_0|redist1|delay_signals[0][105]~q ),
	.ena(en[0]),
	.q(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[20]~q ),
	.prn(vcc));
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[20] .is_wysiwyg = "true";
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[20] .power_up = "low";

dffeas \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[21] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][72]~q ),
	.asdata(\fp_functions_0|redist1|delay_signals[0][73]~q ),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\fp_functions_0|redist1|delay_signals[0][105]~q ),
	.ena(en[0]),
	.q(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[21]~q ),
	.prn(vcc));
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[21] .is_wysiwyg = "true";
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[21] .power_up = "low";

dffeas \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[22] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][73]~q ),
	.asdata(\fp_functions_0|redist1|delay_signals[0][74]~q ),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\fp_functions_0|redist1|delay_signals[0][105]~q ),
	.ena(en[0]),
	.q(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[22]~q ),
	.prn(vcc));
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[22] .is_wysiwyg = "true";
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[22] .power_up = "low";

dffeas \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[23] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][74]~q ),
	.asdata(\fp_functions_0|redist1|delay_signals[0][75]~q ),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\fp_functions_0|redist1|delay_signals[0][105]~q ),
	.ena(en[0]),
	.q(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[23]~q ),
	.prn(vcc));
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[23] .is_wysiwyg = "true";
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[23] .power_up = "low";

dffeas \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[24] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][75]~q ),
	.asdata(\fp_functions_0|redist1|delay_signals[0][76]~q ),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\fp_functions_0|redist1|delay_signals[0][105]~q ),
	.ena(en[0]),
	.q(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[24]~q ),
	.prn(vcc));
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[24] .is_wysiwyg = "true";
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[24] .power_up = "low";

dffeas \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[25] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][76]~q ),
	.asdata(\fp_functions_0|redist1|delay_signals[0][77]~q ),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\fp_functions_0|redist1|delay_signals[0][105]~q ),
	.ena(en[0]),
	.q(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[25]~q ),
	.prn(vcc));
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[25] .is_wysiwyg = "true";
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[25] .power_up = "low";

dffeas \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[26] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][77]~q ),
	.asdata(\fp_functions_0|redist1|delay_signals[0][78]~q ),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\fp_functions_0|redist1|delay_signals[0][105]~q ),
	.ena(en[0]),
	.q(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[26]~q ),
	.prn(vcc));
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[26] .is_wysiwyg = "true";
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[26] .power_up = "low";

dffeas \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[27] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][78]~q ),
	.asdata(\fp_functions_0|redist1|delay_signals[0][79]~q ),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\fp_functions_0|redist1|delay_signals[0][105]~q ),
	.ena(en[0]),
	.q(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[27]~q ),
	.prn(vcc));
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[27] .is_wysiwyg = "true";
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[27] .power_up = "low";

dffeas \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[28] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][79]~q ),
	.asdata(\fp_functions_0|redist1|delay_signals[0][80]~q ),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\fp_functions_0|redist1|delay_signals[0][105]~q ),
	.ena(en[0]),
	.q(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[28]~q ),
	.prn(vcc));
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[28] .is_wysiwyg = "true";
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[28] .power_up = "low";

dffeas \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[29] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][80]~q ),
	.asdata(\fp_functions_0|redist1|delay_signals[0][81]~q ),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\fp_functions_0|redist1|delay_signals[0][105]~q ),
	.ena(en[0]),
	.q(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[29]~q ),
	.prn(vcc));
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[29] .is_wysiwyg = "true";
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[29] .power_up = "low";

dffeas \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[30] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][81]~q ),
	.asdata(\fp_functions_0|redist1|delay_signals[0][82]~q ),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\fp_functions_0|redist1|delay_signals[0][105]~q ),
	.ena(en[0]),
	.q(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[30]~q ),
	.prn(vcc));
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[30] .is_wysiwyg = "true";
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[30] .power_up = "low";

dffeas \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[31] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][82]~q ),
	.asdata(\fp_functions_0|redist1|delay_signals[0][83]~q ),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\fp_functions_0|redist1|delay_signals[0][105]~q ),
	.ena(en[0]),
	.q(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[31]~q ),
	.prn(vcc));
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[31] .is_wysiwyg = "true";
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[31] .power_up = "low";

dffeas \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[32] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][83]~q ),
	.asdata(\fp_functions_0|redist1|delay_signals[0][84]~q ),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\fp_functions_0|redist1|delay_signals[0][105]~q ),
	.ena(en[0]),
	.q(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[32]~q ),
	.prn(vcc));
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[32] .is_wysiwyg = "true";
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[32] .power_up = "low";

dffeas \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[33] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][84]~q ),
	.asdata(\fp_functions_0|redist1|delay_signals[0][85]~q ),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\fp_functions_0|redist1|delay_signals[0][105]~q ),
	.ena(en[0]),
	.q(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[33]~q ),
	.prn(vcc));
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[33] .is_wysiwyg = "true";
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[33] .power_up = "low";

dffeas \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[34] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][85]~q ),
	.asdata(\fp_functions_0|redist1|delay_signals[0][86]~q ),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\fp_functions_0|redist1|delay_signals[0][105]~q ),
	.ena(en[0]),
	.q(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[34]~q ),
	.prn(vcc));
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[34] .is_wysiwyg = "true";
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[34] .power_up = "low";

dffeas \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[35] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][86]~q ),
	.asdata(\fp_functions_0|redist1|delay_signals[0][87]~q ),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\fp_functions_0|redist1|delay_signals[0][105]~q ),
	.ena(en[0]),
	.q(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[35]~q ),
	.prn(vcc));
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[35] .is_wysiwyg = "true";
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[35] .power_up = "low";

dffeas \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[36] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][87]~q ),
	.asdata(\fp_functions_0|redist1|delay_signals[0][88]~q ),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\fp_functions_0|redist1|delay_signals[0][105]~q ),
	.ena(en[0]),
	.q(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[36]~q ),
	.prn(vcc));
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[36] .is_wysiwyg = "true";
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[36] .power_up = "low";

dffeas \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[37] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][88]~q ),
	.asdata(\fp_functions_0|redist1|delay_signals[0][89]~q ),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\fp_functions_0|redist1|delay_signals[0][105]~q ),
	.ena(en[0]),
	.q(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[37]~q ),
	.prn(vcc));
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[37] .is_wysiwyg = "true";
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[37] .power_up = "low";

dffeas \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[38] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][89]~q ),
	.asdata(\fp_functions_0|redist1|delay_signals[0][90]~q ),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\fp_functions_0|redist1|delay_signals[0][105]~q ),
	.ena(en[0]),
	.q(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[38]~q ),
	.prn(vcc));
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[38] .is_wysiwyg = "true";
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[38] .power_up = "low";

dffeas \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[39] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][90]~q ),
	.asdata(\fp_functions_0|redist1|delay_signals[0][91]~q ),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\fp_functions_0|redist1|delay_signals[0][105]~q ),
	.ena(en[0]),
	.q(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[39]~q ),
	.prn(vcc));
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[39] .is_wysiwyg = "true";
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[39] .power_up = "low";

dffeas \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[40] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][91]~q ),
	.asdata(\fp_functions_0|redist1|delay_signals[0][92]~q ),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\fp_functions_0|redist1|delay_signals[0][105]~q ),
	.ena(en[0]),
	.q(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[40]~q ),
	.prn(vcc));
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[40] .is_wysiwyg = "true";
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[40] .power_up = "low";

dffeas \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[41] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][92]~q ),
	.asdata(\fp_functions_0|redist1|delay_signals[0][93]~q ),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\fp_functions_0|redist1|delay_signals[0][105]~q ),
	.ena(en[0]),
	.q(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[41]~q ),
	.prn(vcc));
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[41] .is_wysiwyg = "true";
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[41] .power_up = "low";

dffeas \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[42] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][93]~q ),
	.asdata(\fp_functions_0|redist1|delay_signals[0][94]~q ),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\fp_functions_0|redist1|delay_signals[0][105]~q ),
	.ena(en[0]),
	.q(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[42]~q ),
	.prn(vcc));
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[42] .is_wysiwyg = "true";
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[42] .power_up = "low";

dffeas \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[43] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][94]~q ),
	.asdata(\fp_functions_0|redist1|delay_signals[0][95]~q ),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\fp_functions_0|redist1|delay_signals[0][105]~q ),
	.ena(en[0]),
	.q(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[43]~q ),
	.prn(vcc));
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[43] .is_wysiwyg = "true";
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[43] .power_up = "low";

dffeas \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[44] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][95]~q ),
	.asdata(\fp_functions_0|redist1|delay_signals[0][96]~q ),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\fp_functions_0|redist1|delay_signals[0][105]~q ),
	.ena(en[0]),
	.q(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[44]~q ),
	.prn(vcc));
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[44] .is_wysiwyg = "true";
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[44] .power_up = "low";

dffeas \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[45] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][96]~q ),
	.asdata(\fp_functions_0|redist1|delay_signals[0][97]~q ),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\fp_functions_0|redist1|delay_signals[0][105]~q ),
	.ena(en[0]),
	.q(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[45]~q ),
	.prn(vcc));
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[45] .is_wysiwyg = "true";
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[45] .power_up = "low";

dffeas \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[46] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][97]~q ),
	.asdata(\fp_functions_0|redist1|delay_signals[0][98]~q ),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\fp_functions_0|redist1|delay_signals[0][105]~q ),
	.ena(en[0]),
	.q(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[46]~q ),
	.prn(vcc));
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[46] .is_wysiwyg = "true";
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[46] .power_up = "low";

dffeas \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[47] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][98]~q ),
	.asdata(\fp_functions_0|redist1|delay_signals[0][99]~q ),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\fp_functions_0|redist1|delay_signals[0][105]~q ),
	.ena(en[0]),
	.q(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[47]~q ),
	.prn(vcc));
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[47] .is_wysiwyg = "true";
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[47] .power_up = "low";

dffeas \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[48] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][99]~q ),
	.asdata(\fp_functions_0|redist1|delay_signals[0][100]~q ),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\fp_functions_0|redist1|delay_signals[0][105]~q ),
	.ena(en[0]),
	.q(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[48]~q ),
	.prn(vcc));
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[48] .is_wysiwyg = "true";
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[48] .power_up = "low";

dffeas \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[49] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][100]~q ),
	.asdata(\fp_functions_0|redist1|delay_signals[0][101]~q ),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\fp_functions_0|redist1|delay_signals[0][105]~q ),
	.ena(en[0]),
	.q(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[49]~q ),
	.prn(vcc));
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[49] .is_wysiwyg = "true";
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[49] .power_up = "low";

dffeas \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[50] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][101]~q ),
	.asdata(\fp_functions_0|redist1|delay_signals[0][102]~q ),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\fp_functions_0|redist1|delay_signals[0][105]~q ),
	.ena(en[0]),
	.q(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[50]~q ),
	.prn(vcc));
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[50] .is_wysiwyg = "true";
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[50] .power_up = "low";

dffeas \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[51] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][102]~q ),
	.asdata(\fp_functions_0|redist1|delay_signals[0][103]~q ),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\fp_functions_0|redist1|delay_signals[0][105]~q ),
	.ena(en[0]),
	.q(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[51]~q ),
	.prn(vcc));
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[51] .is_wysiwyg = "true";
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[51] .power_up = "low";

dffeas \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[52] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][103]~q ),
	.asdata(\fp_functions_0|redist1|delay_signals[0][104]~q ),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\fp_functions_0|redist1|delay_signals[0][105]~q ),
	.ena(en[0]),
	.q(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[52]~q ),
	.prn(vcc));
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[52] .is_wysiwyg = "true";
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[52] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|add_5~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist15_outputreg|delay_signals[0][1]~q ),
	.datae(gnd),
	.dataf(!\fp_functions_0|redist15_outputreg|delay_signals[0][0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_5~1_sumout ),
	.cout(\fp_functions_0|add_5~2 ),
	.shareout());
defparam \fp_functions_0|add_5~1 .extended_lut = "off";
defparam \fp_functions_0|add_5~1 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_5~1 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_5~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist15_outputreg|delay_signals[0][2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_5~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_5~5_sumout ),
	.cout(\fp_functions_0|add_5~6 ),
	.shareout());
defparam \fp_functions_0|add_5~5 .extended_lut = "off";
defparam \fp_functions_0|add_5~5 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_5~5 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_5~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist15_outputreg|delay_signals[0][3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_5~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_5~9_sumout ),
	.cout(\fp_functions_0|add_5~10 ),
	.shareout());
defparam \fp_functions_0|add_5~9 .extended_lut = "off";
defparam \fp_functions_0|add_5~9 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_5~9 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_5~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist15_outputreg|delay_signals[0][4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_5~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_5~13_sumout ),
	.cout(\fp_functions_0|add_5~14 ),
	.shareout());
defparam \fp_functions_0|add_5~13 .extended_lut = "off";
defparam \fp_functions_0|add_5~13 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_5~13 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_5~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist15_outputreg|delay_signals[0][5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_5~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_5~17_sumout ),
	.cout(\fp_functions_0|add_5~18 ),
	.shareout());
defparam \fp_functions_0|add_5~17 .extended_lut = "off";
defparam \fp_functions_0|add_5~17 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_5~17 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_5~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist15_outputreg|delay_signals[0][6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_5~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_5~21_sumout ),
	.cout(\fp_functions_0|add_5~22 ),
	.shareout());
defparam \fp_functions_0|add_5~21 .extended_lut = "off";
defparam \fp_functions_0|add_5~21 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_5~21 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_5~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist15_outputreg|delay_signals[0][7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_5~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_5~25_sumout ),
	.cout(\fp_functions_0|add_5~26 ),
	.shareout());
defparam \fp_functions_0|add_5~25 .extended_lut = "off";
defparam \fp_functions_0|add_5~25 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_5~25 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_5~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist15_outputreg|delay_signals[0][8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_5~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_5~29_sumout ),
	.cout(\fp_functions_0|add_5~30 ),
	.shareout());
defparam \fp_functions_0|add_5~29 .extended_lut = "off";
defparam \fp_functions_0|add_5~29 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_5~29 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_5~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist15_outputreg|delay_signals[0][9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_5~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_5~33_sumout ),
	.cout(\fp_functions_0|add_5~34 ),
	.shareout());
defparam \fp_functions_0|add_5~33 .extended_lut = "off";
defparam \fp_functions_0|add_5~33 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_5~33 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_5~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist15_outputreg|delay_signals[0][10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_5~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_5~37_sumout ),
	.cout(\fp_functions_0|add_5~38 ),
	.shareout());
defparam \fp_functions_0|add_5~37 .extended_lut = "off";
defparam \fp_functions_0|add_5~37 .lut_mask = 64'h00000000000000FF;
defparam \fp_functions_0|add_5~37 .shared_arith = "off";

dffeas \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[0] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][51]~q ),
	.asdata(\fp_functions_0|redist1|delay_signals[0][52]~q ),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\fp_functions_0|redist1|delay_signals[0][105]~q ),
	.ena(en[0]),
	.q(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[0]~q ),
	.prn(vcc));
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[0] .is_wysiwyg = "true";
defparam \fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[0] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|add_5~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_5~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_5~41_sumout ),
	.cout(),
	.shareout());
defparam \fp_functions_0|add_5~41 .extended_lut = "off";
defparam \fp_functions_0|add_5~41 .lut_mask = 64'h0000FFFF0000FFFF;
defparam \fp_functions_0|add_5~41 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~265 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][65]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~270 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~265_sumout ),
	.cout(\fp_functions_0|add_6~266 ),
	.shareout());
defparam \fp_functions_0|add_6~265 .extended_lut = "off";
defparam \fp_functions_0|add_6~265 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~265 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_7~18 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist9|delay_signals[0][11]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_7~22_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fp_functions_0|add_7~18_cout ),
	.shareout());
defparam \fp_functions_0|add_7~18 .extended_lut = "off";
defparam \fp_functions_0|add_7~18 .lut_mask = 64'h00000000000000FF;
defparam \fp_functions_0|add_7~18 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_8~18 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist9|delay_signals[0][11]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_8~22_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fp_functions_0|add_8~18_cout ),
	.shareout());
defparam \fp_functions_0|add_8~18 .extended_lut = "off";
defparam \fp_functions_0|add_8~18 .lut_mask = 64'h0000FFFF0000FF00;
defparam \fp_functions_0|add_8~18 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist0|delay_signals[0][27]~q ),
	.datae(gnd),
	.dataf(!\fp_functions_0|redist2|delay_signals[0][27]~q ),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~218 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~1_sumout ),
	.cout(\fp_functions_0|add_1~2 ),
	.shareout());
defparam \fp_functions_0|add_1~1 .extended_lut = "off";
defparam \fp_functions_0|add_1~1 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_1~1 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist0|delay_signals[0][28]~q ),
	.datae(gnd),
	.dataf(!\fp_functions_0|redist2|delay_signals[0][28]~q ),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~5_sumout ),
	.cout(\fp_functions_0|add_1~6 ),
	.shareout());
defparam \fp_functions_0|add_1~5 .extended_lut = "off";
defparam \fp_functions_0|add_1~5 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_1~5 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist2|delay_signals[0][80]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~214 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~9_sumout ),
	.cout(),
	.shareout());
defparam \fp_functions_0|add_1~9 .extended_lut = "off";
defparam \fp_functions_0|add_1~9 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_1~9 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_5~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_5~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_5~45_sumout ),
	.cout(\fp_functions_0|add_5~46 ),
	.shareout());
defparam \fp_functions_0|add_5~45 .extended_lut = "off";
defparam \fp_functions_0|add_5~45 .lut_mask = 64'h0000FFFF0000FFFF;
defparam \fp_functions_0|add_5~45 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_6~269 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist11|delay_signals[0][64]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_6~250 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_6~269_sumout ),
	.cout(\fp_functions_0|add_6~270 ),
	.shareout());
defparam \fp_functions_0|add_6~269 .extended_lut = "off";
defparam \fp_functions_0|add_6~269 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_6~269 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_7~22 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist9|delay_signals[0][10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_7~26_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fp_functions_0|add_7~22_cout ),
	.shareout());
defparam \fp_functions_0|add_7~22 .extended_lut = "off";
defparam \fp_functions_0|add_7~22 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_7~22 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_8~22 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist9|delay_signals[0][10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_8~26_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fp_functions_0|add_8~22_cout ),
	.shareout());
defparam \fp_functions_0|add_8~22 .extended_lut = "off";
defparam \fp_functions_0|add_8~22 .lut_mask = 64'h0000FFFF0000FF00;
defparam \fp_functions_0|add_8~22 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist0|delay_signals[0][29]~q ),
	.datae(gnd),
	.dataf(!\fp_functions_0|redist2|delay_signals[0][29]~q ),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~13_sumout ),
	.cout(\fp_functions_0|add_1~14 ),
	.shareout());
defparam \fp_functions_0|add_1~13 .extended_lut = "off";
defparam \fp_functions_0|add_1~13 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_1~13 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist0|delay_signals[0][30]~q ),
	.datae(gnd),
	.dataf(!\fp_functions_0|redist2|delay_signals[0][30]~q ),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~17_sumout ),
	.cout(\fp_functions_0|add_1~18 ),
	.shareout());
defparam \fp_functions_0|add_1~17 .extended_lut = "off";
defparam \fp_functions_0|add_1~17 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_1~17 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist0|delay_signals[0][31]~q ),
	.datae(gnd),
	.dataf(!\fp_functions_0|redist2|delay_signals[0][31]~q ),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~21_sumout ),
	.cout(\fp_functions_0|add_1~22 ),
	.shareout());
defparam \fp_functions_0|add_1~21 .extended_lut = "off";
defparam \fp_functions_0|add_1~21 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_1~21 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist0|delay_signals[0][32]~q ),
	.datae(gnd),
	.dataf(!\fp_functions_0|redist2|delay_signals[0][32]~q ),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~25_sumout ),
	.cout(\fp_functions_0|add_1~26 ),
	.shareout());
defparam \fp_functions_0|add_1~25 .extended_lut = "off";
defparam \fp_functions_0|add_1~25 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_1~25 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist0|delay_signals[0][33]~q ),
	.datae(gnd),
	.dataf(!\fp_functions_0|redist2|delay_signals[0][33]~q ),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~29_sumout ),
	.cout(\fp_functions_0|add_1~30 ),
	.shareout());
defparam \fp_functions_0|add_1~29 .extended_lut = "off";
defparam \fp_functions_0|add_1~29 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_1~29 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist0|delay_signals[0][34]~q ),
	.datae(gnd),
	.dataf(!\fp_functions_0|redist2|delay_signals[0][34]~q ),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~33_sumout ),
	.cout(\fp_functions_0|add_1~34 ),
	.shareout());
defparam \fp_functions_0|add_1~33 .extended_lut = "off";
defparam \fp_functions_0|add_1~33 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_1~33 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist0|delay_signals[0][35]~q ),
	.datae(gnd),
	.dataf(!\fp_functions_0|redist2|delay_signals[0][35]~q ),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~37_sumout ),
	.cout(\fp_functions_0|add_1~38 ),
	.shareout());
defparam \fp_functions_0|add_1~37 .extended_lut = "off";
defparam \fp_functions_0|add_1~37 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_1~37 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist0|delay_signals[0][36]~q ),
	.datae(gnd),
	.dataf(!\fp_functions_0|redist2|delay_signals[0][36]~q ),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~41_sumout ),
	.cout(\fp_functions_0|add_1~42 ),
	.shareout());
defparam \fp_functions_0|add_1~41 .extended_lut = "off";
defparam \fp_functions_0|add_1~41 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_1~41 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist0|delay_signals[0][37]~q ),
	.datae(gnd),
	.dataf(!\fp_functions_0|redist2|delay_signals[0][37]~q ),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~45_sumout ),
	.cout(\fp_functions_0|add_1~46 ),
	.shareout());
defparam \fp_functions_0|add_1~45 .extended_lut = "off";
defparam \fp_functions_0|add_1~45 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_1~45 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist0|delay_signals[0][38]~q ),
	.datae(gnd),
	.dataf(!\fp_functions_0|redist2|delay_signals[0][38]~q ),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~49_sumout ),
	.cout(\fp_functions_0|add_1~50 ),
	.shareout());
defparam \fp_functions_0|add_1~49 .extended_lut = "off";
defparam \fp_functions_0|add_1~49 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_1~49 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist0|delay_signals[0][39]~q ),
	.datae(gnd),
	.dataf(!\fp_functions_0|redist2|delay_signals[0][39]~q ),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~53_sumout ),
	.cout(\fp_functions_0|add_1~54 ),
	.shareout());
defparam \fp_functions_0|add_1~53 .extended_lut = "off";
defparam \fp_functions_0|add_1~53 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_1~53 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist0|delay_signals[0][40]~q ),
	.datae(gnd),
	.dataf(!\fp_functions_0|redist2|delay_signals[0][40]~q ),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~57_sumout ),
	.cout(\fp_functions_0|add_1~58 ),
	.shareout());
defparam \fp_functions_0|add_1~57 .extended_lut = "off";
defparam \fp_functions_0|add_1~57 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_1~57 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist0|delay_signals[0][41]~q ),
	.datae(gnd),
	.dataf(!\fp_functions_0|redist2|delay_signals[0][41]~q ),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~61_sumout ),
	.cout(\fp_functions_0|add_1~62 ),
	.shareout());
defparam \fp_functions_0|add_1~61 .extended_lut = "off";
defparam \fp_functions_0|add_1~61 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_1~61 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist0|delay_signals[0][42]~q ),
	.datae(gnd),
	.dataf(!\fp_functions_0|redist2|delay_signals[0][42]~q ),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~65_sumout ),
	.cout(\fp_functions_0|add_1~66 ),
	.shareout());
defparam \fp_functions_0|add_1~65 .extended_lut = "off";
defparam \fp_functions_0|add_1~65 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_1~65 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist0|delay_signals[0][43]~q ),
	.datae(gnd),
	.dataf(!\fp_functions_0|redist2|delay_signals[0][43]~q ),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~69_sumout ),
	.cout(\fp_functions_0|add_1~70 ),
	.shareout());
defparam \fp_functions_0|add_1~69 .extended_lut = "off";
defparam \fp_functions_0|add_1~69 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_1~69 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~73 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist0|delay_signals[0][44]~q ),
	.datae(gnd),
	.dataf(!\fp_functions_0|redist2|delay_signals[0][44]~q ),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~73_sumout ),
	.cout(\fp_functions_0|add_1~74 ),
	.shareout());
defparam \fp_functions_0|add_1~73 .extended_lut = "off";
defparam \fp_functions_0|add_1~73 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_1~73 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~77 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist0|delay_signals[0][45]~q ),
	.datae(gnd),
	.dataf(!\fp_functions_0|redist2|delay_signals[0][45]~q ),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~74 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~77_sumout ),
	.cout(\fp_functions_0|add_1~78 ),
	.shareout());
defparam \fp_functions_0|add_1~77 .extended_lut = "off";
defparam \fp_functions_0|add_1~77 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_1~77 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~81 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist0|delay_signals[0][46]~q ),
	.datae(gnd),
	.dataf(!\fp_functions_0|redist2|delay_signals[0][46]~q ),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~78 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~81_sumout ),
	.cout(\fp_functions_0|add_1~82 ),
	.shareout());
defparam \fp_functions_0|add_1~81 .extended_lut = "off";
defparam \fp_functions_0|add_1~81 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_1~81 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~85 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist0|delay_signals[0][47]~q ),
	.datae(gnd),
	.dataf(!\fp_functions_0|redist2|delay_signals[0][47]~q ),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~82 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~85_sumout ),
	.cout(\fp_functions_0|add_1~86 ),
	.shareout());
defparam \fp_functions_0|add_1~85 .extended_lut = "off";
defparam \fp_functions_0|add_1~85 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_1~85 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~89 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist0|delay_signals[0][48]~q ),
	.datae(gnd),
	.dataf(!\fp_functions_0|redist2|delay_signals[0][48]~q ),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~86 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~89_sumout ),
	.cout(\fp_functions_0|add_1~90 ),
	.shareout());
defparam \fp_functions_0|add_1~89 .extended_lut = "off";
defparam \fp_functions_0|add_1~89 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_1~89 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~93 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist0|delay_signals[0][49]~q ),
	.datae(gnd),
	.dataf(!\fp_functions_0|redist2|delay_signals[0][49]~q ),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~90 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~93_sumout ),
	.cout(\fp_functions_0|add_1~94 ),
	.shareout());
defparam \fp_functions_0|add_1~93 .extended_lut = "off";
defparam \fp_functions_0|add_1~93 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_1~93 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~97 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist0|delay_signals[0][50]~q ),
	.datae(gnd),
	.dataf(!\fp_functions_0|redist2|delay_signals[0][50]~q ),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~94 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~97_sumout ),
	.cout(\fp_functions_0|add_1~98 ),
	.shareout());
defparam \fp_functions_0|add_1~97 .extended_lut = "off";
defparam \fp_functions_0|add_1~97 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_1~97 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~101 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist0|delay_signals[0][51]~q ),
	.datae(gnd),
	.dataf(!\fp_functions_0|redist2|delay_signals[0][51]~q ),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~98 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~101_sumout ),
	.cout(\fp_functions_0|add_1~102 ),
	.shareout());
defparam \fp_functions_0|add_1~101 .extended_lut = "off";
defparam \fp_functions_0|add_1~101 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_1~101 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~105 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist0|delay_signals[0][52]~q ),
	.datae(gnd),
	.dataf(!\fp_functions_0|redist2|delay_signals[0][52]~q ),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~102 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~105_sumout ),
	.cout(\fp_functions_0|add_1~106 ),
	.shareout());
defparam \fp_functions_0|add_1~105 .extended_lut = "off";
defparam \fp_functions_0|add_1~105 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_1~105 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~109 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist0|delay_signals[0][53]~q ),
	.datae(gnd),
	.dataf(!\fp_functions_0|redist2|delay_signals[0][53]~q ),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~106 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~109_sumout ),
	.cout(\fp_functions_0|add_1~110 ),
	.shareout());
defparam \fp_functions_0|add_1~109 .extended_lut = "off";
defparam \fp_functions_0|add_1~109 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_1~109 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~113 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist0|delay_signals[0][54]~q ),
	.datae(gnd),
	.dataf(!\fp_functions_0|redist2|delay_signals[0][54]~q ),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~110 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~113_sumout ),
	.cout(\fp_functions_0|add_1~114 ),
	.shareout());
defparam \fp_functions_0|add_1~113 .extended_lut = "off";
defparam \fp_functions_0|add_1~113 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_1~113 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~117 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist2|delay_signals[0][55]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~114 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~117_sumout ),
	.cout(\fp_functions_0|add_1~118 ),
	.shareout());
defparam \fp_functions_0|add_1~117 .extended_lut = "off";
defparam \fp_functions_0|add_1~117 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_1~117 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~121 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist2|delay_signals[0][56]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~118 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~121_sumout ),
	.cout(\fp_functions_0|add_1~122 ),
	.shareout());
defparam \fp_functions_0|add_1~121 .extended_lut = "off";
defparam \fp_functions_0|add_1~121 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_1~121 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~125 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist2|delay_signals[0][57]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~122 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~125_sumout ),
	.cout(\fp_functions_0|add_1~126 ),
	.shareout());
defparam \fp_functions_0|add_1~125 .extended_lut = "off";
defparam \fp_functions_0|add_1~125 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_1~125 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~129 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist2|delay_signals[0][58]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~126 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~129_sumout ),
	.cout(\fp_functions_0|add_1~130 ),
	.shareout());
defparam \fp_functions_0|add_1~129 .extended_lut = "off";
defparam \fp_functions_0|add_1~129 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_1~129 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~133 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist2|delay_signals[0][59]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~130 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~133_sumout ),
	.cout(\fp_functions_0|add_1~134 ),
	.shareout());
defparam \fp_functions_0|add_1~133 .extended_lut = "off";
defparam \fp_functions_0|add_1~133 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_1~133 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~137 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist2|delay_signals[0][60]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~134 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~137_sumout ),
	.cout(\fp_functions_0|add_1~138 ),
	.shareout());
defparam \fp_functions_0|add_1~137 .extended_lut = "off";
defparam \fp_functions_0|add_1~137 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_1~137 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~141 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist2|delay_signals[0][61]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~138 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~141_sumout ),
	.cout(\fp_functions_0|add_1~142 ),
	.shareout());
defparam \fp_functions_0|add_1~141 .extended_lut = "off";
defparam \fp_functions_0|add_1~141 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_1~141 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~145 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist2|delay_signals[0][62]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~142 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~145_sumout ),
	.cout(\fp_functions_0|add_1~146 ),
	.shareout());
defparam \fp_functions_0|add_1~145 .extended_lut = "off";
defparam \fp_functions_0|add_1~145 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_1~145 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~149 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist2|delay_signals[0][63]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~146 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~149_sumout ),
	.cout(\fp_functions_0|add_1~150 ),
	.shareout());
defparam \fp_functions_0|add_1~149 .extended_lut = "off";
defparam \fp_functions_0|add_1~149 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_1~149 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~153 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist2|delay_signals[0][64]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~150 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~153_sumout ),
	.cout(\fp_functions_0|add_1~154 ),
	.shareout());
defparam \fp_functions_0|add_1~153 .extended_lut = "off";
defparam \fp_functions_0|add_1~153 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_1~153 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~157 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist2|delay_signals[0][65]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~154 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~157_sumout ),
	.cout(\fp_functions_0|add_1~158 ),
	.shareout());
defparam \fp_functions_0|add_1~157 .extended_lut = "off";
defparam \fp_functions_0|add_1~157 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_1~157 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~161 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist2|delay_signals[0][66]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~158 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~161_sumout ),
	.cout(\fp_functions_0|add_1~162 ),
	.shareout());
defparam \fp_functions_0|add_1~161 .extended_lut = "off";
defparam \fp_functions_0|add_1~161 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_1~161 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~165 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist2|delay_signals[0][67]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~162 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~165_sumout ),
	.cout(\fp_functions_0|add_1~166 ),
	.shareout());
defparam \fp_functions_0|add_1~165 .extended_lut = "off";
defparam \fp_functions_0|add_1~165 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_1~165 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~169 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist2|delay_signals[0][68]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~166 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~169_sumout ),
	.cout(\fp_functions_0|add_1~170 ),
	.shareout());
defparam \fp_functions_0|add_1~169 .extended_lut = "off";
defparam \fp_functions_0|add_1~169 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_1~169 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~173 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist2|delay_signals[0][69]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~170 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~173_sumout ),
	.cout(\fp_functions_0|add_1~174 ),
	.shareout());
defparam \fp_functions_0|add_1~173 .extended_lut = "off";
defparam \fp_functions_0|add_1~173 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_1~173 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~177 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist2|delay_signals[0][70]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~174 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~177_sumout ),
	.cout(\fp_functions_0|add_1~178 ),
	.shareout());
defparam \fp_functions_0|add_1~177 .extended_lut = "off";
defparam \fp_functions_0|add_1~177 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_1~177 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~181 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist2|delay_signals[0][71]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~178 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~181_sumout ),
	.cout(\fp_functions_0|add_1~182 ),
	.shareout());
defparam \fp_functions_0|add_1~181 .extended_lut = "off";
defparam \fp_functions_0|add_1~181 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_1~181 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~185 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist2|delay_signals[0][72]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~182 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~185_sumout ),
	.cout(\fp_functions_0|add_1~186 ),
	.shareout());
defparam \fp_functions_0|add_1~185 .extended_lut = "off";
defparam \fp_functions_0|add_1~185 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_1~185 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~189 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist2|delay_signals[0][73]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~186 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~189_sumout ),
	.cout(\fp_functions_0|add_1~190 ),
	.shareout());
defparam \fp_functions_0|add_1~189 .extended_lut = "off";
defparam \fp_functions_0|add_1~189 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_1~189 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~193 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist2|delay_signals[0][74]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~190 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~193_sumout ),
	.cout(\fp_functions_0|add_1~194 ),
	.shareout());
defparam \fp_functions_0|add_1~193 .extended_lut = "off";
defparam \fp_functions_0|add_1~193 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_1~193 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~197 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist2|delay_signals[0][75]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~194 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~197_sumout ),
	.cout(\fp_functions_0|add_1~198 ),
	.shareout());
defparam \fp_functions_0|add_1~197 .extended_lut = "off";
defparam \fp_functions_0|add_1~197 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_1~197 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~201 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist2|delay_signals[0][76]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~198 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~201_sumout ),
	.cout(\fp_functions_0|add_1~202 ),
	.shareout());
defparam \fp_functions_0|add_1~201 .extended_lut = "off";
defparam \fp_functions_0|add_1~201 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_1~201 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~205 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist2|delay_signals[0][77]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~202 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~205_sumout ),
	.cout(\fp_functions_0|add_1~206 ),
	.shareout());
defparam \fp_functions_0|add_1~205 .extended_lut = "off";
defparam \fp_functions_0|add_1~205 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_1~205 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~209 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist2|delay_signals[0][78]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~206 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~209_sumout ),
	.cout(\fp_functions_0|add_1~210 ),
	.shareout());
defparam \fp_functions_0|add_1~209 .extended_lut = "off";
defparam \fp_functions_0|add_1~209 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_1~209 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~213 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist2|delay_signals[0][79]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~210 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~213_sumout ),
	.cout(\fp_functions_0|add_1~214 ),
	.shareout());
defparam \fp_functions_0|add_1~213 .extended_lut = "off";
defparam \fp_functions_0|add_1~213 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_1~213 .shared_arith = "off";

twentynm_mlab_cell \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0 (
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.ena2(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\fp_functions_0|redist15_inputreg|delay_signals[0][0]~q }),
	.portaaddr({gnd,gnd,gnd,\fp_functions_0|redist15_wraddr_q[1]~q ,\fp_functions_0|redist15_wraddr_q[0]~q }),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,gnd,\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|rdaddr_reg[1]~q ,\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|rdaddr_reg[0]~q }),
	.portbdataout(\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0_PORTBDATAOUT_bus ));
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0 .address_width = 2;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0 .data_width = 1;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0 .first_address = 0;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0 .first_bit_number = 0;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0 .init_file = "none";
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0 .last_address = 2;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0 .logical_ram_depth = 3;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0 .logical_ram_name = "fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0";
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0 .logical_ram_width = 12;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama0 .mixed_port_feed_through_mode = "dont care";

twentynm_lcell_comb \fp_functions_0|add_1~217 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist0|delay_signals[0][26]~q ),
	.datae(gnd),
	.dataf(!\fp_functions_0|redist2|delay_signals[0][26]~q ),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~230 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~217_sumout ),
	.cout(\fp_functions_0|add_1~218 ),
	.shareout());
defparam \fp_functions_0|add_1~217 .extended_lut = "off";
defparam \fp_functions_0|add_1~217 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_1~217 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~221 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist0|delay_signals[0][23]~q ),
	.datae(gnd),
	.dataf(!\fp_functions_0|redist2|delay_signals[0][23]~q ),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~242 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~221_sumout ),
	.cout(\fp_functions_0|add_1~222 ),
	.shareout());
defparam \fp_functions_0|add_1~221 .extended_lut = "off";
defparam \fp_functions_0|add_1~221 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_1~221 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~225 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist0|delay_signals[0][24]~q ),
	.datae(gnd),
	.dataf(!\fp_functions_0|redist2|delay_signals[0][24]~q ),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~222 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~225_sumout ),
	.cout(\fp_functions_0|add_1~226 ),
	.shareout());
defparam \fp_functions_0|add_1~225 .extended_lut = "off";
defparam \fp_functions_0|add_1~225 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_1~225 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~229 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist0|delay_signals[0][25]~q ),
	.datae(gnd),
	.dataf(!\fp_functions_0|redist2|delay_signals[0][25]~q ),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~226 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~229_sumout ),
	.cout(\fp_functions_0|add_1~230 ),
	.shareout());
defparam \fp_functions_0|add_1~229 .extended_lut = "off";
defparam \fp_functions_0|add_1~229 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_1~229 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~233 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist0|delay_signals[0][16]~q ),
	.datae(gnd),
	.dataf(!\fp_functions_0|redist2|delay_signals[0][16]~q ),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~278 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~233_sumout ),
	.cout(\fp_functions_0|add_1~234 ),
	.shareout());
defparam \fp_functions_0|add_1~233 .extended_lut = "off";
defparam \fp_functions_0|add_1~233 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_1~233 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~237 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist0|delay_signals[0][21]~q ),
	.datae(gnd),
	.dataf(!\fp_functions_0|redist2|delay_signals[0][21]~q ),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~258 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~237_sumout ),
	.cout(\fp_functions_0|add_1~238 ),
	.shareout());
defparam \fp_functions_0|add_1~237 .extended_lut = "off";
defparam \fp_functions_0|add_1~237 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_1~237 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~241 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist0|delay_signals[0][22]~q ),
	.datae(gnd),
	.dataf(!\fp_functions_0|redist2|delay_signals[0][22]~q ),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~238 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~241_sumout ),
	.cout(\fp_functions_0|add_1~242 ),
	.shareout());
defparam \fp_functions_0|add_1~241 .extended_lut = "off";
defparam \fp_functions_0|add_1~241 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_1~241 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~245 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist0|delay_signals[0][17]~q ),
	.datae(gnd),
	.dataf(!\fp_functions_0|redist2|delay_signals[0][17]~q ),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~234 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~245_sumout ),
	.cout(\fp_functions_0|add_1~246 ),
	.shareout());
defparam \fp_functions_0|add_1~245 .extended_lut = "off";
defparam \fp_functions_0|add_1~245 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_1~245 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~249 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist0|delay_signals[0][18]~q ),
	.datae(gnd),
	.dataf(!\fp_functions_0|redist2|delay_signals[0][18]~q ),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~246 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~249_sumout ),
	.cout(\fp_functions_0|add_1~250 ),
	.shareout());
defparam \fp_functions_0|add_1~249 .extended_lut = "off";
defparam \fp_functions_0|add_1~249 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_1~249 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~253 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist0|delay_signals[0][19]~q ),
	.datae(gnd),
	.dataf(!\fp_functions_0|redist2|delay_signals[0][19]~q ),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~250 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~253_sumout ),
	.cout(\fp_functions_0|add_1~254 ),
	.shareout());
defparam \fp_functions_0|add_1~253 .extended_lut = "off";
defparam \fp_functions_0|add_1~253 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_1~253 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~257 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist0|delay_signals[0][20]~q ),
	.datae(gnd),
	.dataf(!\fp_functions_0|redist2|delay_signals[0][20]~q ),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~254 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~257_sumout ),
	.cout(\fp_functions_0|add_1~258 ),
	.shareout());
defparam \fp_functions_0|add_1~257 .extended_lut = "off";
defparam \fp_functions_0|add_1~257 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_1~257 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~261 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist0|delay_signals[0][11]~q ),
	.datae(gnd),
	.dataf(!\fp_functions_0|redist2|delay_signals[0][11]~q ),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~286 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~261_sumout ),
	.cout(\fp_functions_0|add_1~262 ),
	.shareout());
defparam \fp_functions_0|add_1~261 .extended_lut = "off";
defparam \fp_functions_0|add_1~261 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_1~261 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~265 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist0|delay_signals[0][12]~q ),
	.datae(gnd),
	.dataf(!\fp_functions_0|redist2|delay_signals[0][12]~q ),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~262 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~265_sumout ),
	.cout(\fp_functions_0|add_1~266 ),
	.shareout());
defparam \fp_functions_0|add_1~265 .extended_lut = "off";
defparam \fp_functions_0|add_1~265 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_1~265 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~269 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist0|delay_signals[0][13]~q ),
	.datae(gnd),
	.dataf(!\fp_functions_0|redist2|delay_signals[0][13]~q ),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~266 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~269_sumout ),
	.cout(\fp_functions_0|add_1~270 ),
	.shareout());
defparam \fp_functions_0|add_1~269 .extended_lut = "off";
defparam \fp_functions_0|add_1~269 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_1~269 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~273 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist0|delay_signals[0][14]~q ),
	.datae(gnd),
	.dataf(!\fp_functions_0|redist2|delay_signals[0][14]~q ),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~270 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~273_sumout ),
	.cout(\fp_functions_0|add_1~274 ),
	.shareout());
defparam \fp_functions_0|add_1~273 .extended_lut = "off";
defparam \fp_functions_0|add_1~273 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_1~273 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~277 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist0|delay_signals[0][15]~q ),
	.datae(gnd),
	.dataf(!\fp_functions_0|redist2|delay_signals[0][15]~q ),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~274 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~277_sumout ),
	.cout(\fp_functions_0|add_1~278 ),
	.shareout());
defparam \fp_functions_0|add_1~277 .extended_lut = "off";
defparam \fp_functions_0|add_1~277 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_1~277 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~281 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist0|delay_signals[0][4]~q ),
	.datae(gnd),
	.dataf(!\fp_functions_0|redist2|delay_signals[0][4]~q ),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~302 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~281_sumout ),
	.cout(\fp_functions_0|add_1~282 ),
	.shareout());
defparam \fp_functions_0|add_1~281 .extended_lut = "off";
defparam \fp_functions_0|add_1~281 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_1~281 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~285 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist0|delay_signals[0][10]~q ),
	.datae(gnd),
	.dataf(!\fp_functions_0|redist2|delay_signals[0][10]~q ),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~322 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~285_sumout ),
	.cout(\fp_functions_0|add_1~286 ),
	.shareout());
defparam \fp_functions_0|add_1~285 .extended_lut = "off";
defparam \fp_functions_0|add_1~285 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_1~285 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~289 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist0|delay_signals[0][0]~q ),
	.datae(gnd),
	.dataf(!\fp_functions_0|redist2|delay_signals[0][0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~289_sumout ),
	.cout(\fp_functions_0|add_1~290 ),
	.shareout());
defparam \fp_functions_0|add_1~289 .extended_lut = "off";
defparam \fp_functions_0|add_1~289 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_1~289 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~293 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist0|delay_signals[0][1]~q ),
	.datae(gnd),
	.dataf(!\fp_functions_0|redist2|delay_signals[0][1]~q ),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~290 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~293_sumout ),
	.cout(\fp_functions_0|add_1~294 ),
	.shareout());
defparam \fp_functions_0|add_1~293 .extended_lut = "off";
defparam \fp_functions_0|add_1~293 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_1~293 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~297 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist0|delay_signals[0][2]~q ),
	.datae(gnd),
	.dataf(!\fp_functions_0|redist2|delay_signals[0][2]~q ),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~294 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~297_sumout ),
	.cout(\fp_functions_0|add_1~298 ),
	.shareout());
defparam \fp_functions_0|add_1~297 .extended_lut = "off";
defparam \fp_functions_0|add_1~297 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_1~297 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~301 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist0|delay_signals[0][3]~q ),
	.datae(gnd),
	.dataf(!\fp_functions_0|redist2|delay_signals[0][3]~q ),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~298 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~301_sumout ),
	.cout(\fp_functions_0|add_1~302 ),
	.shareout());
defparam \fp_functions_0|add_1~301 .extended_lut = "off";
defparam \fp_functions_0|add_1~301 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_1~301 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~305 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist0|delay_signals[0][5]~q ),
	.datae(gnd),
	.dataf(!\fp_functions_0|redist2|delay_signals[0][5]~q ),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~282 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~305_sumout ),
	.cout(\fp_functions_0|add_1~306 ),
	.shareout());
defparam \fp_functions_0|add_1~305 .extended_lut = "off";
defparam \fp_functions_0|add_1~305 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_1~305 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~309 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist0|delay_signals[0][6]~q ),
	.datae(gnd),
	.dataf(!\fp_functions_0|redist2|delay_signals[0][6]~q ),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~306 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~309_sumout ),
	.cout(\fp_functions_0|add_1~310 ),
	.shareout());
defparam \fp_functions_0|add_1~309 .extended_lut = "off";
defparam \fp_functions_0|add_1~309 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_1~309 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~313 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist0|delay_signals[0][7]~q ),
	.datae(gnd),
	.dataf(!\fp_functions_0|redist2|delay_signals[0][7]~q ),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~310 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~313_sumout ),
	.cout(\fp_functions_0|add_1~314 ),
	.shareout());
defparam \fp_functions_0|add_1~313 .extended_lut = "off";
defparam \fp_functions_0|add_1~313 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_1~313 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~317 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist0|delay_signals[0][8]~q ),
	.datae(gnd),
	.dataf(!\fp_functions_0|redist2|delay_signals[0][8]~q ),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~314 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~317_sumout ),
	.cout(\fp_functions_0|add_1~318 ),
	.shareout());
defparam \fp_functions_0|add_1~317 .extended_lut = "off";
defparam \fp_functions_0|add_1~317 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_1~317 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_1~321 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist0|delay_signals[0][9]~q ),
	.datae(gnd),
	.dataf(!\fp_functions_0|redist2|delay_signals[0][9]~q ),
	.datag(gnd),
	.cin(\fp_functions_0|add_1~318 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_1~321_sumout ),
	.cout(\fp_functions_0|add_1~322 ),
	.shareout());
defparam \fp_functions_0|add_1~321 .extended_lut = "off";
defparam \fp_functions_0|add_1~321 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_1~321 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_5~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist15_outputreg|delay_signals[0][11]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_5~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_5~49_sumout ),
	.cout(\fp_functions_0|add_5~50 ),
	.shareout());
defparam \fp_functions_0|add_5~49 .extended_lut = "off";
defparam \fp_functions_0|add_5~49 .lut_mask = 64'h00000000000000FF;
defparam \fp_functions_0|add_5~49 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_7~26 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist9|delay_signals[0][9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_7~30_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fp_functions_0|add_7~26_cout ),
	.shareout());
defparam \fp_functions_0|add_7~26 .extended_lut = "off";
defparam \fp_functions_0|add_7~26 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_7~26 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_8~26 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist9|delay_signals[0][9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_8~30_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fp_functions_0|add_8~26_cout ),
	.shareout());
defparam \fp_functions_0|add_8~26 .extended_lut = "off";
defparam \fp_functions_0|add_8~26 .lut_mask = 64'h0000FFFF0000FF00;
defparam \fp_functions_0|add_8~26 .shared_arith = "off";

twentynm_mlab_cell \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1 (
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.ena2(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\fp_functions_0|redist15_inputreg|delay_signals[0][1]~q }),
	.portaaddr({gnd,gnd,gnd,\fp_functions_0|redist15_wraddr_q[1]~q ,\fp_functions_0|redist15_wraddr_q[0]~q }),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,gnd,\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|rdaddr_reg[1]~q ,\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|rdaddr_reg[0]~q }),
	.portbdataout(\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1_PORTBDATAOUT_bus ));
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1 .address_width = 2;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1 .data_width = 1;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1 .first_address = 0;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1 .first_bit_number = 1;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1 .init_file = "none";
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1 .last_address = 2;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1 .logical_ram_depth = 3;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1 .logical_ram_name = "fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1";
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1 .logical_ram_width = 12;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama1 .mixed_port_feed_through_mode = "dont care";

twentynm_mlab_cell \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2 (
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.ena2(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\fp_functions_0|redist15_inputreg|delay_signals[0][2]~q }),
	.portaaddr({gnd,gnd,gnd,\fp_functions_0|redist15_wraddr_q[1]~q ,\fp_functions_0|redist15_wraddr_q[0]~q }),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,gnd,\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|rdaddr_reg[1]~q ,\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|rdaddr_reg[0]~q }),
	.portbdataout(\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2_PORTBDATAOUT_bus ));
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2 .address_width = 2;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2 .data_width = 1;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2 .first_address = 0;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2 .first_bit_number = 2;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2 .init_file = "none";
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2 .last_address = 2;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2 .logical_ram_depth = 3;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2 .logical_ram_name = "fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2";
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2 .logical_ram_width = 12;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama2 .mixed_port_feed_through_mode = "dont care";

twentynm_mlab_cell \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3 (
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.ena2(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\fp_functions_0|redist15_inputreg|delay_signals[0][3]~q }),
	.portaaddr({gnd,gnd,gnd,\fp_functions_0|redist15_wraddr_q[1]~q ,\fp_functions_0|redist15_wraddr_q[0]~q }),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,gnd,\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|rdaddr_reg[1]~q ,\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|rdaddr_reg[0]~q }),
	.portbdataout(\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3_PORTBDATAOUT_bus ));
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3 .address_width = 2;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3 .data_width = 1;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3 .first_address = 0;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3 .first_bit_number = 3;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3 .init_file = "none";
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3 .last_address = 2;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3 .logical_ram_depth = 3;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3 .logical_ram_name = "fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3";
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3 .logical_ram_width = 12;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama3 .mixed_port_feed_through_mode = "dont care";

twentynm_mlab_cell \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4 (
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.ena2(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\fp_functions_0|redist15_inputreg|delay_signals[0][4]~q }),
	.portaaddr({gnd,gnd,gnd,\fp_functions_0|redist15_wraddr_q[1]~q ,\fp_functions_0|redist15_wraddr_q[0]~q }),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,gnd,\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|rdaddr_reg[1]~q ,\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|rdaddr_reg[0]~q }),
	.portbdataout(\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4_PORTBDATAOUT_bus ));
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4 .address_width = 2;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4 .data_width = 1;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4 .first_address = 0;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4 .first_bit_number = 4;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4 .init_file = "none";
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4 .last_address = 2;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4 .logical_ram_depth = 3;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4 .logical_ram_name = "fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4";
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4 .logical_ram_width = 12;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama4 .mixed_port_feed_through_mode = "dont care";

twentynm_mlab_cell \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5 (
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.ena2(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\fp_functions_0|redist15_inputreg|delay_signals[0][5]~q }),
	.portaaddr({gnd,gnd,gnd,\fp_functions_0|redist15_wraddr_q[1]~q ,\fp_functions_0|redist15_wraddr_q[0]~q }),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,gnd,\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|rdaddr_reg[1]~q ,\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|rdaddr_reg[0]~q }),
	.portbdataout(\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5_PORTBDATAOUT_bus ));
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5 .address_width = 2;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5 .data_width = 1;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5 .first_address = 0;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5 .first_bit_number = 5;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5 .init_file = "none";
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5 .last_address = 2;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5 .logical_ram_depth = 3;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5 .logical_ram_name = "fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5";
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5 .logical_ram_width = 12;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama5 .mixed_port_feed_through_mode = "dont care";

twentynm_mlab_cell \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6 (
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.ena2(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\fp_functions_0|redist15_inputreg|delay_signals[0][6]~q }),
	.portaaddr({gnd,gnd,gnd,\fp_functions_0|redist15_wraddr_q[1]~q ,\fp_functions_0|redist15_wraddr_q[0]~q }),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,gnd,\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|rdaddr_reg[1]~q ,\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|rdaddr_reg[0]~q }),
	.portbdataout(\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6_PORTBDATAOUT_bus ));
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6 .address_width = 2;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6 .data_width = 1;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6 .first_address = 0;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6 .first_bit_number = 6;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6 .init_file = "none";
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6 .last_address = 2;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6 .logical_ram_depth = 3;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6 .logical_ram_name = "fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6";
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6 .logical_ram_width = 12;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama6 .mixed_port_feed_through_mode = "dont care";

twentynm_mlab_cell \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7 (
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.ena2(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\fp_functions_0|redist15_inputreg|delay_signals[0][7]~q }),
	.portaaddr({gnd,gnd,gnd,\fp_functions_0|redist15_wraddr_q[1]~q ,\fp_functions_0|redist15_wraddr_q[0]~q }),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,gnd,\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|rdaddr_reg[1]~q ,\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|rdaddr_reg[0]~q }),
	.portbdataout(\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7_PORTBDATAOUT_bus ));
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7 .address_width = 2;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7 .data_width = 1;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7 .first_address = 0;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7 .first_bit_number = 7;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7 .init_file = "none";
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7 .last_address = 2;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7 .logical_ram_depth = 3;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7 .logical_ram_name = "fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7";
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7 .logical_ram_width = 12;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama7 .mixed_port_feed_through_mode = "dont care";

twentynm_mlab_cell \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8 (
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.ena2(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\fp_functions_0|redist15_inputreg|delay_signals[0][8]~q }),
	.portaaddr({gnd,gnd,gnd,\fp_functions_0|redist15_wraddr_q[1]~q ,\fp_functions_0|redist15_wraddr_q[0]~q }),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,gnd,\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|rdaddr_reg[1]~q ,\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|rdaddr_reg[0]~q }),
	.portbdataout(\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8_PORTBDATAOUT_bus ));
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8 .address_width = 2;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8 .data_width = 1;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8 .first_address = 0;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8 .first_bit_number = 8;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8 .init_file = "none";
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8 .last_address = 2;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8 .logical_ram_depth = 3;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8 .logical_ram_name = "fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8";
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8 .logical_ram_width = 12;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama8 .mixed_port_feed_through_mode = "dont care";

twentynm_mlab_cell \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9 (
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.ena2(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\fp_functions_0|redist15_inputreg|delay_signals[0][9]~q }),
	.portaaddr({gnd,gnd,gnd,\fp_functions_0|redist15_wraddr_q[1]~q ,\fp_functions_0|redist15_wraddr_q[0]~q }),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,gnd,\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|rdaddr_reg[1]~q ,\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|rdaddr_reg[0]~q }),
	.portbdataout(\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9_PORTBDATAOUT_bus ));
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9 .address_width = 2;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9 .data_width = 1;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9 .first_address = 0;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9 .first_bit_number = 9;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9 .init_file = "none";
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9 .last_address = 2;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9 .logical_ram_depth = 3;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9 .logical_ram_name = "fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9";
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9 .logical_ram_width = 12;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama9 .mixed_port_feed_through_mode = "dont care";

twentynm_mlab_cell \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10 (
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.ena2(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\fp_functions_0|redist15_inputreg|delay_signals[0][10]~q }),
	.portaaddr({gnd,gnd,gnd,\fp_functions_0|redist15_wraddr_q[1]~q ,\fp_functions_0|redist15_wraddr_q[0]~q }),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,gnd,\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|rdaddr_reg[1]~q ,\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|rdaddr_reg[0]~q }),
	.portbdataout(\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10_PORTBDATAOUT_bus ));
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10 .address_width = 2;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10 .data_width = 1;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10 .first_address = 0;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10 .first_bit_number = 10;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10 .init_file = "none";
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10 .last_address = 2;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10 .logical_ram_depth = 3;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10 .logical_ram_name = "fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10";
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10 .logical_ram_width = 12;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama10 .mixed_port_feed_through_mode = "dont care";

twentynm_lcell_comb \fp_functions_0|add_7~30 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist9|delay_signals[0][8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_7~34_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fp_functions_0|add_7~30_cout ),
	.shareout());
defparam \fp_functions_0|add_7~30 .extended_lut = "off";
defparam \fp_functions_0|add_7~30 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_7~30 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_8~30 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist9|delay_signals[0][8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_8~34_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fp_functions_0|add_8~30_cout ),
	.shareout());
defparam \fp_functions_0|add_8~30 .extended_lut = "off";
defparam \fp_functions_0|add_8~30 .lut_mask = 64'h0000FFFF0000FF00;
defparam \fp_functions_0|add_8~30 .shared_arith = "off";

twentynm_mac \fp_functions_0|mult_2~mac (
	.sub(gnd),
	.negate(gnd),
	.accumulate(gnd),
	.loadconst(gnd),
	.ax({\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][26]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][25]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][24]~q ,
\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][23]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][22]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][21]~q ,
\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][20]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][19]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][18]~q ,
\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][17]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][16]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][15]~q ,
\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][14]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][13]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][12]~q ,
\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][11]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][10]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][9]~q ,
\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][8]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][7]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][6]~q ,
\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][5]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][4]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][3]~q ,
\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][2]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][1]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][0]~q }),
	.ay({\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][26]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][25]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][24]~q ,
\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][23]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][22]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][21]~q ,
\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][20]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][19]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][18]~q ,
\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][17]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][16]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][15]~q ,
\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][14]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][13]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][12]~q ,
\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][11]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][10]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][9]~q ,
\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][8]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][7]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][6]~q ,
\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][5]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][4]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][3]~q ,
\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][2]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][1]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][0]~q }),
	.az(26'b00000000000000000000000000),
	.bx(18'b000000000000000000),
	.by(19'b0000000000000000000),
	.bz(18'b000000000000000000),
	.coefsela(3'b000),
	.coefselb(3'b000),
	.clk(3'b000),
	.aclr(2'b00),
	.ena(3'b111),
	.scanin(27'b000000000000000000000000000),
	.chainin({\fp_functions_0|mult_3~149 ,\fp_functions_0|mult_3~148 ,\fp_functions_0|mult_3~147 ,\fp_functions_0|mult_3~146 ,\fp_functions_0|mult_3~145 ,\fp_functions_0|mult_3~144 ,\fp_functions_0|mult_3~143 ,\fp_functions_0|mult_3~142 ,\fp_functions_0|mult_3~141 ,
\fp_functions_0|mult_3~140 ,\fp_functions_0|mult_3~139 ,\fp_functions_0|mult_3~138 ,\fp_functions_0|mult_3~137 ,\fp_functions_0|mult_3~136 ,\fp_functions_0|mult_3~135 ,\fp_functions_0|mult_3~134 ,\fp_functions_0|mult_3~133 ,\fp_functions_0|mult_3~132 ,
\fp_functions_0|mult_3~131 ,\fp_functions_0|mult_3~130 ,\fp_functions_0|mult_3~129 ,\fp_functions_0|mult_3~128 ,\fp_functions_0|mult_3~127 ,\fp_functions_0|mult_3~126 ,\fp_functions_0|mult_3~125 ,\fp_functions_0|mult_3~124 ,\fp_functions_0|mult_3~123 ,
\fp_functions_0|mult_3~122 ,\fp_functions_0|mult_3~121 ,\fp_functions_0|mult_3~120 ,\fp_functions_0|mult_3~119 ,\fp_functions_0|mult_3~118 ,\fp_functions_0|mult_3~117 ,\fp_functions_0|mult_3~116 ,\fp_functions_0|mult_3~115 ,\fp_functions_0|mult_3~114 ,
\fp_functions_0|mult_3~113 ,\fp_functions_0|mult_3~112 ,\fp_functions_0|mult_3~111 ,\fp_functions_0|mult_3~110 ,\fp_functions_0|mult_3~109 ,\fp_functions_0|mult_3~108 ,\fp_functions_0|mult_3~107 ,\fp_functions_0|mult_3~106 ,\fp_functions_0|mult_3~105 ,
\fp_functions_0|mult_3~104 ,\fp_functions_0|mult_3~103 ,\fp_functions_0|mult_3~102 ,\fp_functions_0|mult_3~101 ,\fp_functions_0|mult_3~100 ,\fp_functions_0|mult_3~99 ,\fp_functions_0|mult_3~98 ,\fp_functions_0|mult_3~97 ,\fp_functions_0|mult_3~96 ,
\fp_functions_0|mult_3~95 ,\fp_functions_0|mult_3~94 ,\fp_functions_0|mult_3~93 ,\fp_functions_0|mult_3~92 ,\fp_functions_0|mult_3~91 ,\fp_functions_0|mult_3~90 ,\fp_functions_0|mult_3~89 ,\fp_functions_0|mult_3~88 ,\fp_functions_0|mult_3~87 ,
\fp_functions_0|mult_3~86 }),
	.dftout(),
	.resulta(\fp_functions_0|mult_2~mac_RESULTA_bus ),
	.resultb(),
	.scanout(),
	.chainout());
defparam \fp_functions_0|mult_2~mac .accum_pipeline_clock = "none";
defparam \fp_functions_0|mult_2~mac .accumulate_clock = "none";
defparam \fp_functions_0|mult_2~mac .ax_clock = "none";
defparam \fp_functions_0|mult_2~mac .ax_width = 27;
defparam \fp_functions_0|mult_2~mac .ay_scan_in_clock = "none";
defparam \fp_functions_0|mult_2~mac .ay_scan_in_width = 27;
defparam \fp_functions_0|mult_2~mac .ay_use_scan_in = "false";
defparam \fp_functions_0|mult_2~mac .az_clock = "none";
defparam \fp_functions_0|mult_2~mac .bx_clock = "none";
defparam \fp_functions_0|mult_2~mac .by_clock = "none";
defparam \fp_functions_0|mult_2~mac .by_use_scan_in = "false";
defparam \fp_functions_0|mult_2~mac .bz_clock = "none";
defparam \fp_functions_0|mult_2~mac .coef_a_0 = 0;
defparam \fp_functions_0|mult_2~mac .coef_a_1 = 0;
defparam \fp_functions_0|mult_2~mac .coef_a_2 = 0;
defparam \fp_functions_0|mult_2~mac .coef_a_3 = 0;
defparam \fp_functions_0|mult_2~mac .coef_a_4 = 0;
defparam \fp_functions_0|mult_2~mac .coef_a_5 = 0;
defparam \fp_functions_0|mult_2~mac .coef_a_6 = 0;
defparam \fp_functions_0|mult_2~mac .coef_a_7 = 0;
defparam \fp_functions_0|mult_2~mac .coef_b_0 = 0;
defparam \fp_functions_0|mult_2~mac .coef_b_1 = 0;
defparam \fp_functions_0|mult_2~mac .coef_b_2 = 0;
defparam \fp_functions_0|mult_2~mac .coef_b_3 = 0;
defparam \fp_functions_0|mult_2~mac .coef_b_4 = 0;
defparam \fp_functions_0|mult_2~mac .coef_b_5 = 0;
defparam \fp_functions_0|mult_2~mac .coef_b_6 = 0;
defparam \fp_functions_0|mult_2~mac .coef_b_7 = 0;
defparam \fp_functions_0|mult_2~mac .coef_sel_a_clock = "none";
defparam \fp_functions_0|mult_2~mac .coef_sel_b_clock = "none";
defparam \fp_functions_0|mult_2~mac .delay_scan_out_ay = "false";
defparam \fp_functions_0|mult_2~mac .delay_scan_out_by = "false";
defparam \fp_functions_0|mult_2~mac .enable_double_accum = "false";
defparam \fp_functions_0|mult_2~mac .input_pipeline_clock = "none";
defparam \fp_functions_0|mult_2~mac .load_const_clock = "none";
defparam \fp_functions_0|mult_2~mac .load_const_pipeline_clock = "none";
defparam \fp_functions_0|mult_2~mac .load_const_value = 0;
defparam \fp_functions_0|mult_2~mac .mode_sub_location = 0;
defparam \fp_functions_0|mult_2~mac .negate_clock = "none";
defparam \fp_functions_0|mult_2~mac .negate_pipeline_clock = "none";
defparam \fp_functions_0|mult_2~mac .operand_source_max = "input";
defparam \fp_functions_0|mult_2~mac .operand_source_may = "input";
defparam \fp_functions_0|mult_2~mac .operand_source_mbx = "input";
defparam \fp_functions_0|mult_2~mac .operand_source_mby = "input";
defparam \fp_functions_0|mult_2~mac .operation_mode = "m27x27";
defparam \fp_functions_0|mult_2~mac .output_clock = "none";
defparam \fp_functions_0|mult_2~mac .preadder_subtract_a = "false";
defparam \fp_functions_0|mult_2~mac .preadder_subtract_b = "false";
defparam \fp_functions_0|mult_2~mac .result_a_width = 64;
defparam \fp_functions_0|mult_2~mac .signed_max = "false";
defparam \fp_functions_0|mult_2~mac .signed_may = "false";
defparam \fp_functions_0|mult_2~mac .signed_mbx = "false";
defparam \fp_functions_0|mult_2~mac .signed_mby = "false";
defparam \fp_functions_0|mult_2~mac .sub_clock = "none";
defparam \fp_functions_0|mult_2~mac .sub_pipeline_clock = "none";
defparam \fp_functions_0|mult_2~mac .use_chainadder = "true";

twentynm_mac \fp_functions_0|mult_0~mac (
	.sub(gnd),
	.negate(gnd),
	.accumulate(gnd),
	.loadconst(gnd),
	.ax({\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][26]~q ,\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][25]~q ,\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][24]~q ,
\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][23]~q ,\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][22]~q ,\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][21]~q ,
\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][20]~q ,\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][19]~q ,\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][18]~q ,
\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][17]~q ,\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][16]~q ,\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][15]~q ,
\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][14]~q ,\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][13]~q ,\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][12]~q ,
\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][11]~q ,\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][10]~q ,\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][9]~q ,
\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][8]~q ,\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][7]~q ,\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][6]~q ,
\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][5]~q ,\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][4]~q ,\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][3]~q ,
\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][2]~q ,\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][1]~q ,\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][0]~q }),
	.ay({\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][26]~q ,\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][25]~q ,\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][24]~q ,
\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][23]~q ,\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][22]~q ,\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][21]~q ,
\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][20]~q ,\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][19]~q ,\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][18]~q ,
\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][17]~q ,\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][16]~q ,\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][15]~q ,
\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][14]~q ,\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][13]~q ,\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][12]~q ,
\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][11]~q ,\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][10]~q ,\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][9]~q ,
\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][8]~q ,\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][7]~q ,\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][6]~q ,
\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][5]~q ,\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][4]~q ,\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][3]~q ,
\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][2]~q ,\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][1]~q ,\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][0]~q }),
	.az(26'b00000000000000000000000000),
	.bx(18'b000000000000000000),
	.by(19'b0000000000000000000),
	.bz(18'b000000000000000000),
	.coefsela(3'b000),
	.coefselb(3'b000),
	.clk(3'b000),
	.aclr(2'b00),
	.ena(3'b111),
	.scanin(27'b000000000000000000000000000),
	.chainin(1'b0),
	.dftout(),
	.resulta(\fp_functions_0|mult_0~mac_RESULTA_bus ),
	.resultb(),
	.scanout(),
	.chainout());
defparam \fp_functions_0|mult_0~mac .accum_pipeline_clock = "none";
defparam \fp_functions_0|mult_0~mac .accumulate_clock = "none";
defparam \fp_functions_0|mult_0~mac .ax_clock = "none";
defparam \fp_functions_0|mult_0~mac .ax_width = 27;
defparam \fp_functions_0|mult_0~mac .ay_scan_in_clock = "none";
defparam \fp_functions_0|mult_0~mac .ay_scan_in_width = 27;
defparam \fp_functions_0|mult_0~mac .ay_use_scan_in = "false";
defparam \fp_functions_0|mult_0~mac .az_clock = "none";
defparam \fp_functions_0|mult_0~mac .bx_clock = "none";
defparam \fp_functions_0|mult_0~mac .by_clock = "none";
defparam \fp_functions_0|mult_0~mac .by_use_scan_in = "false";
defparam \fp_functions_0|mult_0~mac .bz_clock = "none";
defparam \fp_functions_0|mult_0~mac .coef_a_0 = 0;
defparam \fp_functions_0|mult_0~mac .coef_a_1 = 0;
defparam \fp_functions_0|mult_0~mac .coef_a_2 = 0;
defparam \fp_functions_0|mult_0~mac .coef_a_3 = 0;
defparam \fp_functions_0|mult_0~mac .coef_a_4 = 0;
defparam \fp_functions_0|mult_0~mac .coef_a_5 = 0;
defparam \fp_functions_0|mult_0~mac .coef_a_6 = 0;
defparam \fp_functions_0|mult_0~mac .coef_a_7 = 0;
defparam \fp_functions_0|mult_0~mac .coef_b_0 = 0;
defparam \fp_functions_0|mult_0~mac .coef_b_1 = 0;
defparam \fp_functions_0|mult_0~mac .coef_b_2 = 0;
defparam \fp_functions_0|mult_0~mac .coef_b_3 = 0;
defparam \fp_functions_0|mult_0~mac .coef_b_4 = 0;
defparam \fp_functions_0|mult_0~mac .coef_b_5 = 0;
defparam \fp_functions_0|mult_0~mac .coef_b_6 = 0;
defparam \fp_functions_0|mult_0~mac .coef_b_7 = 0;
defparam \fp_functions_0|mult_0~mac .coef_sel_a_clock = "none";
defparam \fp_functions_0|mult_0~mac .coef_sel_b_clock = "none";
defparam \fp_functions_0|mult_0~mac .delay_scan_out_ay = "false";
defparam \fp_functions_0|mult_0~mac .delay_scan_out_by = "false";
defparam \fp_functions_0|mult_0~mac .enable_double_accum = "false";
defparam \fp_functions_0|mult_0~mac .input_pipeline_clock = "none";
defparam \fp_functions_0|mult_0~mac .load_const_clock = "none";
defparam \fp_functions_0|mult_0~mac .load_const_pipeline_clock = "none";
defparam \fp_functions_0|mult_0~mac .load_const_value = 0;
defparam \fp_functions_0|mult_0~mac .mode_sub_location = 0;
defparam \fp_functions_0|mult_0~mac .negate_clock = "none";
defparam \fp_functions_0|mult_0~mac .negate_pipeline_clock = "none";
defparam \fp_functions_0|mult_0~mac .operand_source_max = "input";
defparam \fp_functions_0|mult_0~mac .operand_source_may = "input";
defparam \fp_functions_0|mult_0~mac .operand_source_mbx = "input";
defparam \fp_functions_0|mult_0~mac .operand_source_mby = "input";
defparam \fp_functions_0|mult_0~mac .operation_mode = "m27x27";
defparam \fp_functions_0|mult_0~mac .output_clock = "none";
defparam \fp_functions_0|mult_0~mac .preadder_subtract_a = "false";
defparam \fp_functions_0|mult_0~mac .preadder_subtract_b = "false";
defparam \fp_functions_0|mult_0~mac .result_a_width = 64;
defparam \fp_functions_0|mult_0~mac .signed_max = "false";
defparam \fp_functions_0|mult_0~mac .signed_may = "false";
defparam \fp_functions_0|mult_0~mac .signed_mbx = "false";
defparam \fp_functions_0|mult_0~mac .signed_mby = "false";
defparam \fp_functions_0|mult_0~mac .sub_clock = "none";
defparam \fp_functions_0|mult_0~mac .sub_pipeline_clock = "none";
defparam \fp_functions_0|mult_0~mac .use_chainadder = "false";

twentynm_mac \fp_functions_0|mult_1~12 (
	.sub(gnd),
	.negate(gnd),
	.accumulate(gnd),
	.loadconst(gnd),
	.ax({\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][26]~q ,\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][25]~q ,\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][24]~q ,\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][23]~q ,
\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][22]~q ,\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][21]~q ,\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][20]~q ,\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][19]~q ,
\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][18]~q ,\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][17]~q ,\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][16]~q ,\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][15]~q ,
\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][14]~q ,\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][13]~q ,\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][12]~q ,\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][11]~q ,
\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][10]~q ,\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][9]~q ,\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][8]~q ,\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][7]~q ,
\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][6]~q ,\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][5]~q ,\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][4]~q ,\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][3]~q ,
\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][2]~q ,\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][1]~q ,\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][0]~q }),
	.ay({\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][26]~q ,\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][25]~q ,\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][24]~q ,\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][23]~q ,
\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][22]~q ,\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][21]~q ,\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][20]~q ,\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][19]~q ,
\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][18]~q ,\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][17]~q ,\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][16]~q ,\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][15]~q ,
\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][14]~q ,\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][13]~q ,\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][12]~q ,\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][11]~q ,
\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][10]~q ,\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][9]~q ,\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][8]~q ,\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][7]~q ,
\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][6]~q ,\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][5]~q ,\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][4]~q ,\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][3]~q ,
\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][2]~q ,\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][1]~q ,\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][0]~q }),
	.az(26'b00000000000000000000000000),
	.bx(18'b000000000000000000),
	.by(19'b0000000000000000000),
	.bz(18'b000000000000000000),
	.coefsela(3'b000),
	.coefselb(3'b000),
	.clk(3'b000),
	.aclr(2'b00),
	.ena(3'b111),
	.scanin(27'b000000000000000000000000000),
	.chainin(1'b0),
	.dftout(),
	.resulta(\fp_functions_0|mult_1~12_RESULTA_bus ),
	.resultb(),
	.scanout(),
	.chainout());
defparam \fp_functions_0|mult_1~12 .accum_pipeline_clock = "none";
defparam \fp_functions_0|mult_1~12 .accumulate_clock = "none";
defparam \fp_functions_0|mult_1~12 .ax_clock = "none";
defparam \fp_functions_0|mult_1~12 .ax_width = 27;
defparam \fp_functions_0|mult_1~12 .ay_scan_in_clock = "none";
defparam \fp_functions_0|mult_1~12 .ay_scan_in_width = 27;
defparam \fp_functions_0|mult_1~12 .ay_use_scan_in = "false";
defparam \fp_functions_0|mult_1~12 .az_clock = "none";
defparam \fp_functions_0|mult_1~12 .bx_clock = "none";
defparam \fp_functions_0|mult_1~12 .by_clock = "none";
defparam \fp_functions_0|mult_1~12 .by_use_scan_in = "false";
defparam \fp_functions_0|mult_1~12 .bz_clock = "none";
defparam \fp_functions_0|mult_1~12 .coef_a_0 = 0;
defparam \fp_functions_0|mult_1~12 .coef_a_1 = 0;
defparam \fp_functions_0|mult_1~12 .coef_a_2 = 0;
defparam \fp_functions_0|mult_1~12 .coef_a_3 = 0;
defparam \fp_functions_0|mult_1~12 .coef_a_4 = 0;
defparam \fp_functions_0|mult_1~12 .coef_a_5 = 0;
defparam \fp_functions_0|mult_1~12 .coef_a_6 = 0;
defparam \fp_functions_0|mult_1~12 .coef_a_7 = 0;
defparam \fp_functions_0|mult_1~12 .coef_b_0 = 0;
defparam \fp_functions_0|mult_1~12 .coef_b_1 = 0;
defparam \fp_functions_0|mult_1~12 .coef_b_2 = 0;
defparam \fp_functions_0|mult_1~12 .coef_b_3 = 0;
defparam \fp_functions_0|mult_1~12 .coef_b_4 = 0;
defparam \fp_functions_0|mult_1~12 .coef_b_5 = 0;
defparam \fp_functions_0|mult_1~12 .coef_b_6 = 0;
defparam \fp_functions_0|mult_1~12 .coef_b_7 = 0;
defparam \fp_functions_0|mult_1~12 .coef_sel_a_clock = "none";
defparam \fp_functions_0|mult_1~12 .coef_sel_b_clock = "none";
defparam \fp_functions_0|mult_1~12 .delay_scan_out_ay = "false";
defparam \fp_functions_0|mult_1~12 .delay_scan_out_by = "false";
defparam \fp_functions_0|mult_1~12 .enable_double_accum = "false";
defparam \fp_functions_0|mult_1~12 .input_pipeline_clock = "none";
defparam \fp_functions_0|mult_1~12 .load_const_clock = "none";
defparam \fp_functions_0|mult_1~12 .load_const_pipeline_clock = "none";
defparam \fp_functions_0|mult_1~12 .load_const_value = 0;
defparam \fp_functions_0|mult_1~12 .mode_sub_location = 0;
defparam \fp_functions_0|mult_1~12 .negate_clock = "none";
defparam \fp_functions_0|mult_1~12 .negate_pipeline_clock = "none";
defparam \fp_functions_0|mult_1~12 .operand_source_max = "input";
defparam \fp_functions_0|mult_1~12 .operand_source_may = "input";
defparam \fp_functions_0|mult_1~12 .operand_source_mbx = "input";
defparam \fp_functions_0|mult_1~12 .operand_source_mby = "input";
defparam \fp_functions_0|mult_1~12 .operation_mode = "m27x27";
defparam \fp_functions_0|mult_1~12 .output_clock = "none";
defparam \fp_functions_0|mult_1~12 .preadder_subtract_a = "false";
defparam \fp_functions_0|mult_1~12 .preadder_subtract_b = "false";
defparam \fp_functions_0|mult_1~12 .result_a_width = 64;
defparam \fp_functions_0|mult_1~12 .signed_max = "false";
defparam \fp_functions_0|mult_1~12 .signed_may = "false";
defparam \fp_functions_0|mult_1~12 .signed_mbx = "false";
defparam \fp_functions_0|mult_1~12 .signed_mby = "false";
defparam \fp_functions_0|mult_1~12 .sub_clock = "none";
defparam \fp_functions_0|mult_1~12 .sub_pipeline_clock = "none";
defparam \fp_functions_0|mult_1~12 .use_chainadder = "false";

twentynm_lcell_comb \fp_functions_0|add_7~34 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist9|delay_signals[0][7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_7~38_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fp_functions_0|add_7~34_cout ),
	.shareout());
defparam \fp_functions_0|add_7~34 .extended_lut = "off";
defparam \fp_functions_0|add_7~34 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_7~34 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_8~34 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist9|delay_signals[0][7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_8~38_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fp_functions_0|add_8~34_cout ),
	.shareout());
defparam \fp_functions_0|add_8~34 .extended_lut = "off";
defparam \fp_functions_0|add_8~34 .lut_mask = 64'h0000FFFF0000FF00;
defparam \fp_functions_0|add_8~34 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_4~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!b[52]),
	.datae(gnd),
	.dataf(!a[52]),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_4~1_sumout ),
	.cout(\fp_functions_0|add_4~2 ),
	.shareout());
defparam \fp_functions_0|add_4~1 .extended_lut = "off";
defparam \fp_functions_0|add_4~1 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_4~1 .shared_arith = "off";

twentynm_mac \fp_functions_0|mult_3~mac (
	.sub(gnd),
	.negate(gnd),
	.accumulate(gnd),
	.loadconst(gnd),
	.ax({\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][26]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][25]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][24]~q ,
\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][23]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][22]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][21]~q ,
\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][20]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][19]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][18]~q ,
\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][17]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][16]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][15]~q ,
\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][14]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][13]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][12]~q ,
\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][11]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][10]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][9]~q ,
\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][8]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][7]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][6]~q ,
\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][5]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][4]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][3]~q ,
\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][2]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][1]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][0]~q }),
	.ay({\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][26]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][25]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][24]~q ,
\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][23]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][22]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][21]~q ,
\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][20]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][19]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][18]~q ,
\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][17]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][16]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][15]~q ,
\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][14]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][13]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][12]~q ,
\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][11]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][10]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][9]~q ,
\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][8]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][7]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][6]~q ,
\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][5]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][4]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][3]~q ,
\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][2]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][1]~q ,\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][0]~q }),
	.az(26'b00000000000000000000000000),
	.bx(18'b000000000000000000),
	.by(19'b0000000000000000000),
	.bz(18'b000000000000000000),
	.coefsela(3'b000),
	.coefselb(3'b000),
	.clk({gnd,gnd,clk}),
	.aclr({areset,gnd}),
	.ena({gnd,gnd,en[0]}),
	.scanin(27'b000000000000000000000000000),
	.chainin(1'b0),
	.dftout(),
	.resulta(\fp_functions_0|mult_3~mac_RESULTA_bus ),
	.resultb(),
	.scanout(),
	.chainout(\fp_functions_0|mult_3~mac_CHAINOUT_bus ));
defparam \fp_functions_0|mult_3~mac .accum_pipeline_clock = "none";
defparam \fp_functions_0|mult_3~mac .accumulate_clock = "none";
defparam \fp_functions_0|mult_3~mac .ax_clock = "none";
defparam \fp_functions_0|mult_3~mac .ax_width = 27;
defparam \fp_functions_0|mult_3~mac .ay_scan_in_clock = "none";
defparam \fp_functions_0|mult_3~mac .ay_scan_in_width = 27;
defparam \fp_functions_0|mult_3~mac .ay_use_scan_in = "false";
defparam \fp_functions_0|mult_3~mac .az_clock = "none";
defparam \fp_functions_0|mult_3~mac .bx_clock = "none";
defparam \fp_functions_0|mult_3~mac .by_clock = "none";
defparam \fp_functions_0|mult_3~mac .by_use_scan_in = "false";
defparam \fp_functions_0|mult_3~mac .bz_clock = "none";
defparam \fp_functions_0|mult_3~mac .coef_a_0 = 0;
defparam \fp_functions_0|mult_3~mac .coef_a_1 = 0;
defparam \fp_functions_0|mult_3~mac .coef_a_2 = 0;
defparam \fp_functions_0|mult_3~mac .coef_a_3 = 0;
defparam \fp_functions_0|mult_3~mac .coef_a_4 = 0;
defparam \fp_functions_0|mult_3~mac .coef_a_5 = 0;
defparam \fp_functions_0|mult_3~mac .coef_a_6 = 0;
defparam \fp_functions_0|mult_3~mac .coef_a_7 = 0;
defparam \fp_functions_0|mult_3~mac .coef_b_0 = 0;
defparam \fp_functions_0|mult_3~mac .coef_b_1 = 0;
defparam \fp_functions_0|mult_3~mac .coef_b_2 = 0;
defparam \fp_functions_0|mult_3~mac .coef_b_3 = 0;
defparam \fp_functions_0|mult_3~mac .coef_b_4 = 0;
defparam \fp_functions_0|mult_3~mac .coef_b_5 = 0;
defparam \fp_functions_0|mult_3~mac .coef_b_6 = 0;
defparam \fp_functions_0|mult_3~mac .coef_b_7 = 0;
defparam \fp_functions_0|mult_3~mac .coef_sel_a_clock = "none";
defparam \fp_functions_0|mult_3~mac .coef_sel_b_clock = "none";
defparam \fp_functions_0|mult_3~mac .delay_scan_out_ay = "false";
defparam \fp_functions_0|mult_3~mac .delay_scan_out_by = "false";
defparam \fp_functions_0|mult_3~mac .enable_double_accum = "false";
defparam \fp_functions_0|mult_3~mac .input_pipeline_clock = "none";
defparam \fp_functions_0|mult_3~mac .load_const_clock = "none";
defparam \fp_functions_0|mult_3~mac .load_const_pipeline_clock = "none";
defparam \fp_functions_0|mult_3~mac .load_const_value = 0;
defparam \fp_functions_0|mult_3~mac .mode_sub_location = 0;
defparam \fp_functions_0|mult_3~mac .negate_clock = "none";
defparam \fp_functions_0|mult_3~mac .negate_pipeline_clock = "none";
defparam \fp_functions_0|mult_3~mac .operand_source_max = "input";
defparam \fp_functions_0|mult_3~mac .operand_source_may = "input";
defparam \fp_functions_0|mult_3~mac .operand_source_mbx = "input";
defparam \fp_functions_0|mult_3~mac .operand_source_mby = "input";
defparam \fp_functions_0|mult_3~mac .operation_mode = "m27x27";
defparam \fp_functions_0|mult_3~mac .output_clock = "0";
defparam \fp_functions_0|mult_3~mac .preadder_subtract_a = "false";
defparam \fp_functions_0|mult_3~mac .preadder_subtract_b = "false";
defparam \fp_functions_0|mult_3~mac .result_a_width = 64;
defparam \fp_functions_0|mult_3~mac .signed_max = "false";
defparam \fp_functions_0|mult_3~mac .signed_may = "false";
defparam \fp_functions_0|mult_3~mac .signed_mbx = "false";
defparam \fp_functions_0|mult_3~mac .signed_mby = "false";
defparam \fp_functions_0|mult_3~mac .sub_clock = "none";
defparam \fp_functions_0|mult_3~mac .sub_pipeline_clock = "none";
defparam \fp_functions_0|mult_3~mac .use_chainadder = "false";

twentynm_mlab_cell \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11 (
	.clk0(clk),
	.clk1(gnd),
	.ena0(en[0]),
	.ena1(vcc),
	.ena2(vcc),
	.clr(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\fp_functions_0|redist15_inputreg|delay_signals[0][11]~q }),
	.portaaddr({gnd,gnd,gnd,\fp_functions_0|redist15_wraddr_q[1]~q ,\fp_functions_0|redist15_wraddr_q[0]~q }),
	.portabyteenamasks(1'b1),
	.portbaddr({gnd,gnd,gnd,\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|rdaddr_reg[1]~q ,\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|rdaddr_reg[0]~q }),
	.portbdataout(\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11_PORTBDATAOUT_bus ));
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11 .address_width = 2;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11 .data_width = 1;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11 .first_address = 0;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11 .first_bit_number = 11;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11 .init_file = "none";
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11 .last_address = 2;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11 .logical_ram_depth = 3;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11 .logical_ram_name = "fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11";
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11 .logical_ram_width = 12;
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|lutrama11 .mixed_port_feed_through_mode = "dont care";

twentynm_lcell_comb \fp_functions_0|add_7~38 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist9|delay_signals[0][6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_7~42_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fp_functions_0|add_7~38_cout ),
	.shareout());
defparam \fp_functions_0|add_7~38 .extended_lut = "off";
defparam \fp_functions_0|add_7~38 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_7~38 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_8~38 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist9|delay_signals[0][6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_8~42_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fp_functions_0|add_8~38_cout ),
	.shareout());
defparam \fp_functions_0|add_8~38 .extended_lut = "off";
defparam \fp_functions_0|add_8~38 .lut_mask = 64'h0000FFFF0000FF00;
defparam \fp_functions_0|add_8~38 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_4~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!b[53]),
	.datae(gnd),
	.dataf(!a[53]),
	.datag(gnd),
	.cin(\fp_functions_0|add_4~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_4~5_sumout ),
	.cout(\fp_functions_0|add_4~6 ),
	.shareout());
defparam \fp_functions_0|add_4~5 .extended_lut = "off";
defparam \fp_functions_0|add_4~5 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_4~5 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_4~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!b[54]),
	.datae(gnd),
	.dataf(!a[54]),
	.datag(gnd),
	.cin(\fp_functions_0|add_4~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_4~9_sumout ),
	.cout(\fp_functions_0|add_4~10 ),
	.shareout());
defparam \fp_functions_0|add_4~9 .extended_lut = "off";
defparam \fp_functions_0|add_4~9 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_4~9 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_4~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!b[55]),
	.datae(gnd),
	.dataf(!a[55]),
	.datag(gnd),
	.cin(\fp_functions_0|add_4~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_4~13_sumout ),
	.cout(\fp_functions_0|add_4~14 ),
	.shareout());
defparam \fp_functions_0|add_4~13 .extended_lut = "off";
defparam \fp_functions_0|add_4~13 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_4~13 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_4~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!b[56]),
	.datae(gnd),
	.dataf(!a[56]),
	.datag(gnd),
	.cin(\fp_functions_0|add_4~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_4~17_sumout ),
	.cout(\fp_functions_0|add_4~18 ),
	.shareout());
defparam \fp_functions_0|add_4~17 .extended_lut = "off";
defparam \fp_functions_0|add_4~17 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_4~17 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_4~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!b[57]),
	.datae(gnd),
	.dataf(!a[57]),
	.datag(gnd),
	.cin(\fp_functions_0|add_4~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_4~21_sumout ),
	.cout(\fp_functions_0|add_4~22 ),
	.shareout());
defparam \fp_functions_0|add_4~21 .extended_lut = "off";
defparam \fp_functions_0|add_4~21 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_4~21 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_4~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!b[58]),
	.datae(gnd),
	.dataf(!a[58]),
	.datag(gnd),
	.cin(\fp_functions_0|add_4~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_4~25_sumout ),
	.cout(\fp_functions_0|add_4~26 ),
	.shareout());
defparam \fp_functions_0|add_4~25 .extended_lut = "off";
defparam \fp_functions_0|add_4~25 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_4~25 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_4~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!b[59]),
	.datae(gnd),
	.dataf(!a[59]),
	.datag(gnd),
	.cin(\fp_functions_0|add_4~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_4~29_sumout ),
	.cout(\fp_functions_0|add_4~30 ),
	.shareout());
defparam \fp_functions_0|add_4~29 .extended_lut = "off";
defparam \fp_functions_0|add_4~29 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_4~29 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_4~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!b[60]),
	.datae(gnd),
	.dataf(!a[60]),
	.datag(gnd),
	.cin(\fp_functions_0|add_4~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_4~33_sumout ),
	.cout(\fp_functions_0|add_4~34 ),
	.shareout());
defparam \fp_functions_0|add_4~33 .extended_lut = "off";
defparam \fp_functions_0|add_4~33 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_4~33 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_4~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!b[61]),
	.datae(gnd),
	.dataf(!a[61]),
	.datag(gnd),
	.cin(\fp_functions_0|add_4~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_4~37_sumout ),
	.cout(\fp_functions_0|add_4~38 ),
	.shareout());
defparam \fp_functions_0|add_4~37 .extended_lut = "off";
defparam \fp_functions_0|add_4~37 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_4~37 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_4~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!b[62]),
	.datae(gnd),
	.dataf(!a[62]),
	.datag(gnd),
	.cin(\fp_functions_0|add_4~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_4~41_sumout ),
	.cout(\fp_functions_0|add_4~42 ),
	.shareout());
defparam \fp_functions_0|add_4~41 .extended_lut = "off";
defparam \fp_functions_0|add_4~41 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_4~41 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_7~42 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist9|delay_signals[0][5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_7~46_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fp_functions_0|add_7~42_cout ),
	.shareout());
defparam \fp_functions_0|add_7~42 .extended_lut = "off";
defparam \fp_functions_0|add_7~42 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_7~42 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_8~42 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist9|delay_signals[0][5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_8~46_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fp_functions_0|add_8~42_cout ),
	.shareout());
defparam \fp_functions_0|add_8~42 .extended_lut = "off";
defparam \fp_functions_0|add_8~42 .lut_mask = 64'h0000FFFF0000FF00;
defparam \fp_functions_0|add_8~42 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_7~46 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist9|delay_signals[0][4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_7~50_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fp_functions_0|add_7~46_cout ),
	.shareout());
defparam \fp_functions_0|add_7~46 .extended_lut = "off";
defparam \fp_functions_0|add_7~46 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_7~46 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_8~46 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist9|delay_signals[0][4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_8~50_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fp_functions_0|add_8~46_cout ),
	.shareout());
defparam \fp_functions_0|add_8~46 .extended_lut = "off";
defparam \fp_functions_0|add_8~46 .lut_mask = 64'h0000FFFF0000FF00;
defparam \fp_functions_0|add_8~46 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_4~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_4~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\fp_functions_0|add_4~45_sumout ),
	.cout(),
	.shareout());
defparam \fp_functions_0|add_4~45 .extended_lut = "off";
defparam \fp_functions_0|add_4~45 .lut_mask = 64'h0000FFFF00000000;
defparam \fp_functions_0|add_4~45 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_7~50 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist9|delay_signals[0][3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_7~54_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fp_functions_0|add_7~50_cout ),
	.shareout());
defparam \fp_functions_0|add_7~50 .extended_lut = "off";
defparam \fp_functions_0|add_7~50 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_7~50 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_8~50 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist9|delay_signals[0][3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_8~54_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fp_functions_0|add_8~50_cout ),
	.shareout());
defparam \fp_functions_0|add_8~50 .extended_lut = "off";
defparam \fp_functions_0|add_8~50 .lut_mask = 64'h0000FFFF0000FF00;
defparam \fp_functions_0|add_8~50 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_7~54 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist9|delay_signals[0][2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_7~58_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fp_functions_0|add_7~54_cout ),
	.shareout());
defparam \fp_functions_0|add_7~54 .extended_lut = "off";
defparam \fp_functions_0|add_7~54 .lut_mask = 64'h0000FFFF000000FF;
defparam \fp_functions_0|add_7~54 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_8~54 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist9|delay_signals[0][2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\fp_functions_0|add_8~58_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fp_functions_0|add_8~54_cout ),
	.shareout());
defparam \fp_functions_0|add_8~54 .extended_lut = "off";
defparam \fp_functions_0|add_8~54 .lut_mask = 64'h0000FFFF0000FF00;
defparam \fp_functions_0|add_8~54 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_7~58 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist9|delay_signals[0][1]~q ),
	.datae(gnd),
	.dataf(!\fp_functions_0|redist9|delay_signals[0][0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fp_functions_0|add_7~58_cout ),
	.shareout());
defparam \fp_functions_0|add_7~58 .extended_lut = "off";
defparam \fp_functions_0|add_7~58 .lut_mask = 64'h0000FF00000000FF;
defparam \fp_functions_0|add_7~58 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|add_8~58 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\fp_functions_0|redist9|delay_signals[0][1]~q ),
	.datae(gnd),
	.dataf(!\fp_functions_0|redist9|delay_signals[0][0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\fp_functions_0|add_8~58_cout ),
	.shareout());
defparam \fp_functions_0|add_8~58 .extended_lut = "off";
defparam \fp_functions_0|add_8~58 .lut_mask = 64'h000000FF0000FF00;
defparam \fp_functions_0|add_8~58 .shared_arith = "off";

dffeas \fp_functions_0|redist10|delay_signals[0][0] (
	.clk(clk),
	.d(\fp_functions_0|redist10|delay_signals[1][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[0][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[0][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[0][0] .power_up = "low";

dffeas \fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0] (
	.clk(clk),
	.d(\fp_functions_0|i933~0_combout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0] .is_wysiwyg = "true";
defparam \fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0] .power_up = "low";

dffeas \fp_functions_0|ExcROvfAndInReg_uid84_fpMulTest_delay|delay_signals[0][0] (
	.clk(clk),
	.d(\fp_functions_0|i6384~combout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|ExcROvfAndInReg_uid84_fpMulTest_delay|delay_signals[0][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|ExcROvfAndInReg_uid84_fpMulTest_delay|delay_signals[0][0] .is_wysiwyg = "true";
defparam \fp_functions_0|ExcROvfAndInReg_uid84_fpMulTest_delay|delay_signals[0][0] .power_up = "low";

dffeas \fp_functions_0|excYRAndExcXI_uid83_fpMulTest_delay|delay_signals[0][0] (
	.clk(clk),
	.d(\fp_functions_0|i6387~0_combout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|excYRAndExcXI_uid83_fpMulTest_delay|delay_signals[0][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|excYRAndExcXI_uid83_fpMulTest_delay|delay_signals[0][0] .is_wysiwyg = "true";
defparam \fp_functions_0|excYRAndExcXI_uid83_fpMulTest_delay|delay_signals[0][0] .power_up = "low";

dffeas \fp_functions_0|excXRAndExcYI_uid82_fpMulTest_delay|delay_signals[0][0] (
	.clk(clk),
	.d(\fp_functions_0|i6390~0_combout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|excXRAndExcYI_uid82_fpMulTest_delay|delay_signals[0][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|excXRAndExcYI_uid82_fpMulTest_delay|delay_signals[0][0] .is_wysiwyg = "true";
defparam \fp_functions_0|excXRAndExcYI_uid82_fpMulTest_delay|delay_signals[0][0] .power_up = "low";

dffeas \fp_functions_0|excXIAndExcYI_uid81_fpMulTest_delay|delay_signals[0][0] (
	.clk(clk),
	.d(\fp_functions_0|i6393~0_combout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|excXIAndExcYI_uid81_fpMulTest_delay|delay_signals[0][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|excXIAndExcYI_uid81_fpMulTest_delay|delay_signals[0][0] .is_wysiwyg = "true";
defparam \fp_functions_0|excXIAndExcYI_uid81_fpMulTest_delay|delay_signals[0][0] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|i6400 (
	.dataa(!\fp_functions_0|ExcROvfAndInReg_uid84_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|excYRAndExcXI_uid83_fpMulTest_delay|delay_signals[0][0]~q ),
	.datac(!\fp_functions_0|excXRAndExcYI_uid82_fpMulTest_delay|delay_signals[0][0]~q ),
	.datad(!\fp_functions_0|excXIAndExcYI_uid81_fpMulTest_delay|delay_signals[0][0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|i6400~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|i6400 .extended_lut = "off";
defparam \fp_functions_0|i6400 .lut_mask = 64'h8000800080008000;
defparam \fp_functions_0|i6400 .shared_arith = "off";

dffeas \fp_functions_0|excZC3_uid79_fpMulTest_delay|delay_signals[0][0] (
	.clk(clk),
	.d(\fp_functions_0|i6459~combout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|excZC3_uid79_fpMulTest_delay|delay_signals[0][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|excZC3_uid79_fpMulTest_delay|delay_signals[0][0] .is_wysiwyg = "true";
defparam \fp_functions_0|excZC3_uid79_fpMulTest_delay|delay_signals[0][0] .power_up = "low";

dffeas \fp_functions_0|excYZAndExcXR_uid78_fpMulTest_delay|delay_signals[0][0] (
	.clk(clk),
	.d(\fp_functions_0|i6462~0_combout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|excYZAndExcXR_uid78_fpMulTest_delay|delay_signals[0][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|excYZAndExcXR_uid78_fpMulTest_delay|delay_signals[0][0] .is_wysiwyg = "true";
defparam \fp_functions_0|excYZAndExcXR_uid78_fpMulTest_delay|delay_signals[0][0] .power_up = "low";

dffeas \fp_functions_0|excXZAndExcYR_uid77_fpMulTest_delay|delay_signals[0][0] (
	.clk(clk),
	.d(\fp_functions_0|i6465~0_combout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|excXZAndExcYR_uid77_fpMulTest_delay|delay_signals[0][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|excXZAndExcYR_uid77_fpMulTest_delay|delay_signals[0][0] .is_wysiwyg = "true";
defparam \fp_functions_0|excXZAndExcYR_uid77_fpMulTest_delay|delay_signals[0][0] .power_up = "low";

dffeas \fp_functions_0|excXZAndExcYZ_uid76_fpMulTest_delay|delay_signals[0][0] (
	.clk(clk),
	.d(\fp_functions_0|i6468~combout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|excXZAndExcYZ_uid76_fpMulTest_delay|delay_signals[0][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|excXZAndExcYZ_uid76_fpMulTest_delay|delay_signals[0][0] .is_wysiwyg = "true";
defparam \fp_functions_0|excXZAndExcYZ_uid76_fpMulTest_delay|delay_signals[0][0] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|i6475 (
	.dataa(!\fp_functions_0|excZC3_uid79_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|excYZAndExcXR_uid78_fpMulTest_delay|delay_signals[0][0]~q ),
	.datac(!\fp_functions_0|excXZAndExcYR_uid77_fpMulTest_delay|delay_signals[0][0]~q ),
	.datad(!\fp_functions_0|excXZAndExcYZ_uid76_fpMulTest_delay|delay_signals[0][0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|i6475~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|i6475 .extended_lut = "off";
defparam \fp_functions_0|i6475 .lut_mask = 64'h8000800080008000;
defparam \fp_functions_0|i6475 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|Mux_64~0 (
	.dataa(!\fp_functions_0|redist10|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_64~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_64~0 .extended_lut = "off";
defparam \fp_functions_0|Mux_64~0 .lut_mask = 64'h0007000700070007;
defparam \fp_functions_0|Mux_64~0 .shared_arith = "off";

dffeas \fp_functions_0|redist10|delay_signals[0][1] (
	.clk(clk),
	.d(\fp_functions_0|redist10|delay_signals[1][1]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[0][1]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[0][1] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[0][1] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_63~0 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist10|delay_signals[0][1]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_63~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_63~0 .extended_lut = "off";
defparam \fp_functions_0|Mux_63~0 .lut_mask = 64'h0002000200020002;
defparam \fp_functions_0|Mux_63~0 .shared_arith = "off";

dffeas \fp_functions_0|redist10|delay_signals[0][2] (
	.clk(clk),
	.d(\fp_functions_0|redist10|delay_signals[1][2]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[0][2]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[0][2] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[0][2] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_62~0 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist10|delay_signals[0][2]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_62~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_62~0 .extended_lut = "off";
defparam \fp_functions_0|Mux_62~0 .lut_mask = 64'h0002000200020002;
defparam \fp_functions_0|Mux_62~0 .shared_arith = "off";

dffeas \fp_functions_0|redist10|delay_signals[0][3] (
	.clk(clk),
	.d(\fp_functions_0|redist10|delay_signals[1][3]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[0][3]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[0][3] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[0][3] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_61~0 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist10|delay_signals[0][3]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_61~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_61~0 .extended_lut = "off";
defparam \fp_functions_0|Mux_61~0 .lut_mask = 64'h0002000200020002;
defparam \fp_functions_0|Mux_61~0 .shared_arith = "off";

dffeas \fp_functions_0|redist10|delay_signals[0][4] (
	.clk(clk),
	.d(\fp_functions_0|redist10|delay_signals[1][4]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[0][4]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[0][4] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[0][4] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_60~0 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist10|delay_signals[0][4]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_60~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_60~0 .extended_lut = "off";
defparam \fp_functions_0|Mux_60~0 .lut_mask = 64'h0002000200020002;
defparam \fp_functions_0|Mux_60~0 .shared_arith = "off";

dffeas \fp_functions_0|redist10|delay_signals[0][5] (
	.clk(clk),
	.d(\fp_functions_0|redist10|delay_signals[1][5]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[0][5]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[0][5] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[0][5] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_59~0 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist10|delay_signals[0][5]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_59~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_59~0 .extended_lut = "off";
defparam \fp_functions_0|Mux_59~0 .lut_mask = 64'h0002000200020002;
defparam \fp_functions_0|Mux_59~0 .shared_arith = "off";

dffeas \fp_functions_0|redist10|delay_signals[0][6] (
	.clk(clk),
	.d(\fp_functions_0|redist10|delay_signals[1][6]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[0][6]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[0][6] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[0][6] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_58~0 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist10|delay_signals[0][6]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_58~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_58~0 .extended_lut = "off";
defparam \fp_functions_0|Mux_58~0 .lut_mask = 64'h0002000200020002;
defparam \fp_functions_0|Mux_58~0 .shared_arith = "off";

dffeas \fp_functions_0|redist10|delay_signals[0][7] (
	.clk(clk),
	.d(\fp_functions_0|redist10|delay_signals[1][7]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[0][7]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[0][7] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[0][7] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_57~0 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist10|delay_signals[0][7]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_57~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_57~0 .extended_lut = "off";
defparam \fp_functions_0|Mux_57~0 .lut_mask = 64'h0002000200020002;
defparam \fp_functions_0|Mux_57~0 .shared_arith = "off";

dffeas \fp_functions_0|redist10|delay_signals[0][8] (
	.clk(clk),
	.d(\fp_functions_0|redist10|delay_signals[1][8]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[0][8]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[0][8] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[0][8] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_56~0 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist10|delay_signals[0][8]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_56~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_56~0 .extended_lut = "off";
defparam \fp_functions_0|Mux_56~0 .lut_mask = 64'h0002000200020002;
defparam \fp_functions_0|Mux_56~0 .shared_arith = "off";

dffeas \fp_functions_0|redist10|delay_signals[0][9] (
	.clk(clk),
	.d(\fp_functions_0|redist10|delay_signals[1][9]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[0][9]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[0][9] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[0][9] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_55~0 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist10|delay_signals[0][9]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_55~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_55~0 .extended_lut = "off";
defparam \fp_functions_0|Mux_55~0 .lut_mask = 64'h0002000200020002;
defparam \fp_functions_0|Mux_55~0 .shared_arith = "off";

dffeas \fp_functions_0|redist10|delay_signals[0][10] (
	.clk(clk),
	.d(\fp_functions_0|redist10|delay_signals[1][10]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[0][10]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[0][10] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[0][10] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_54~0 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist10|delay_signals[0][10]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_54~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_54~0 .extended_lut = "off";
defparam \fp_functions_0|Mux_54~0 .lut_mask = 64'h0002000200020002;
defparam \fp_functions_0|Mux_54~0 .shared_arith = "off";

dffeas \fp_functions_0|redist10|delay_signals[0][11] (
	.clk(clk),
	.d(\fp_functions_0|redist10|delay_signals[1][11]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[0][11]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[0][11] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[0][11] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_53~0 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist10|delay_signals[0][11]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_53~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_53~0 .extended_lut = "off";
defparam \fp_functions_0|Mux_53~0 .lut_mask = 64'h0002000200020002;
defparam \fp_functions_0|Mux_53~0 .shared_arith = "off";

dffeas \fp_functions_0|redist10|delay_signals[0][12] (
	.clk(clk),
	.d(\fp_functions_0|redist10|delay_signals[1][12]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[0][12]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[0][12] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[0][12] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_52~0 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist10|delay_signals[0][12]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_52~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_52~0 .extended_lut = "off";
defparam \fp_functions_0|Mux_52~0 .lut_mask = 64'h0002000200020002;
defparam \fp_functions_0|Mux_52~0 .shared_arith = "off";

dffeas \fp_functions_0|redist10|delay_signals[0][13] (
	.clk(clk),
	.d(\fp_functions_0|redist10|delay_signals[1][13]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[0][13]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[0][13] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[0][13] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_51~0 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist10|delay_signals[0][13]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_51~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_51~0 .extended_lut = "off";
defparam \fp_functions_0|Mux_51~0 .lut_mask = 64'h0002000200020002;
defparam \fp_functions_0|Mux_51~0 .shared_arith = "off";

dffeas \fp_functions_0|redist10|delay_signals[0][14] (
	.clk(clk),
	.d(\fp_functions_0|redist10|delay_signals[1][14]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[0][14]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[0][14] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[0][14] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_50~0 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist10|delay_signals[0][14]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_50~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_50~0 .extended_lut = "off";
defparam \fp_functions_0|Mux_50~0 .lut_mask = 64'h0002000200020002;
defparam \fp_functions_0|Mux_50~0 .shared_arith = "off";

dffeas \fp_functions_0|redist10|delay_signals[0][15] (
	.clk(clk),
	.d(\fp_functions_0|redist10|delay_signals[1][15]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[0][15]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[0][15] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[0][15] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_49~0 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist10|delay_signals[0][15]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_49~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_49~0 .extended_lut = "off";
defparam \fp_functions_0|Mux_49~0 .lut_mask = 64'h0002000200020002;
defparam \fp_functions_0|Mux_49~0 .shared_arith = "off";

dffeas \fp_functions_0|redist10|delay_signals[0][16] (
	.clk(clk),
	.d(\fp_functions_0|redist10|delay_signals[1][16]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[0][16]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[0][16] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[0][16] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_48~0 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist10|delay_signals[0][16]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_48~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_48~0 .extended_lut = "off";
defparam \fp_functions_0|Mux_48~0 .lut_mask = 64'h0002000200020002;
defparam \fp_functions_0|Mux_48~0 .shared_arith = "off";

dffeas \fp_functions_0|redist10|delay_signals[0][17] (
	.clk(clk),
	.d(\fp_functions_0|redist10|delay_signals[1][17]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[0][17]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[0][17] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[0][17] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_47~0 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist10|delay_signals[0][17]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_47~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_47~0 .extended_lut = "off";
defparam \fp_functions_0|Mux_47~0 .lut_mask = 64'h0002000200020002;
defparam \fp_functions_0|Mux_47~0 .shared_arith = "off";

dffeas \fp_functions_0|redist10|delay_signals[0][18] (
	.clk(clk),
	.d(\fp_functions_0|redist10|delay_signals[1][18]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[0][18]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[0][18] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[0][18] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_46~0 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist10|delay_signals[0][18]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_46~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_46~0 .extended_lut = "off";
defparam \fp_functions_0|Mux_46~0 .lut_mask = 64'h0002000200020002;
defparam \fp_functions_0|Mux_46~0 .shared_arith = "off";

dffeas \fp_functions_0|redist10|delay_signals[0][19] (
	.clk(clk),
	.d(\fp_functions_0|redist10|delay_signals[1][19]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[0][19]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[0][19] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[0][19] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_45~0 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist10|delay_signals[0][19]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_45~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_45~0 .extended_lut = "off";
defparam \fp_functions_0|Mux_45~0 .lut_mask = 64'h0002000200020002;
defparam \fp_functions_0|Mux_45~0 .shared_arith = "off";

dffeas \fp_functions_0|redist10|delay_signals[0][20] (
	.clk(clk),
	.d(\fp_functions_0|redist10|delay_signals[1][20]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[0][20]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[0][20] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[0][20] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_44~0 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist10|delay_signals[0][20]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_44~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_44~0 .extended_lut = "off";
defparam \fp_functions_0|Mux_44~0 .lut_mask = 64'h0002000200020002;
defparam \fp_functions_0|Mux_44~0 .shared_arith = "off";

dffeas \fp_functions_0|redist10|delay_signals[0][21] (
	.clk(clk),
	.d(\fp_functions_0|redist10|delay_signals[1][21]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[0][21]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[0][21] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[0][21] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_43~0 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist10|delay_signals[0][21]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_43~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_43~0 .extended_lut = "off";
defparam \fp_functions_0|Mux_43~0 .lut_mask = 64'h0002000200020002;
defparam \fp_functions_0|Mux_43~0 .shared_arith = "off";

dffeas \fp_functions_0|redist10|delay_signals[0][22] (
	.clk(clk),
	.d(\fp_functions_0|redist10|delay_signals[1][22]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[0][22]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[0][22] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[0][22] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_42~0 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist10|delay_signals[0][22]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_42~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_42~0 .extended_lut = "off";
defparam \fp_functions_0|Mux_42~0 .lut_mask = 64'h0002000200020002;
defparam \fp_functions_0|Mux_42~0 .shared_arith = "off";

dffeas \fp_functions_0|redist10|delay_signals[0][23] (
	.clk(clk),
	.d(\fp_functions_0|redist10|delay_signals[1][23]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[0][23]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[0][23] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[0][23] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_41~0 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist10|delay_signals[0][23]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_41~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_41~0 .extended_lut = "off";
defparam \fp_functions_0|Mux_41~0 .lut_mask = 64'h0002000200020002;
defparam \fp_functions_0|Mux_41~0 .shared_arith = "off";

dffeas \fp_functions_0|redist10|delay_signals[0][24] (
	.clk(clk),
	.d(\fp_functions_0|redist10|delay_signals[1][24]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[0][24]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[0][24] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[0][24] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_40~0 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist10|delay_signals[0][24]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_40~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_40~0 .extended_lut = "off";
defparam \fp_functions_0|Mux_40~0 .lut_mask = 64'h0002000200020002;
defparam \fp_functions_0|Mux_40~0 .shared_arith = "off";

dffeas \fp_functions_0|redist10|delay_signals[0][25] (
	.clk(clk),
	.d(\fp_functions_0|redist10|delay_signals[1][25]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[0][25]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[0][25] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[0][25] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_39~0 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist10|delay_signals[0][25]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_39~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_39~0 .extended_lut = "off";
defparam \fp_functions_0|Mux_39~0 .lut_mask = 64'h0002000200020002;
defparam \fp_functions_0|Mux_39~0 .shared_arith = "off";

dffeas \fp_functions_0|redist10|delay_signals[0][26] (
	.clk(clk),
	.d(\fp_functions_0|redist10|delay_signals[1][26]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[0][26]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[0][26] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[0][26] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_38~0 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist10|delay_signals[0][26]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_38~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_38~0 .extended_lut = "off";
defparam \fp_functions_0|Mux_38~0 .lut_mask = 64'h0002000200020002;
defparam \fp_functions_0|Mux_38~0 .shared_arith = "off";

dffeas \fp_functions_0|redist10|delay_signals[0][27] (
	.clk(clk),
	.d(\fp_functions_0|redist10|delay_signals[1][27]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[0][27]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[0][27] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[0][27] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_37~0 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist10|delay_signals[0][27]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_37~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_37~0 .extended_lut = "off";
defparam \fp_functions_0|Mux_37~0 .lut_mask = 64'h0002000200020002;
defparam \fp_functions_0|Mux_37~0 .shared_arith = "off";

dffeas \fp_functions_0|redist10|delay_signals[0][28] (
	.clk(clk),
	.d(\fp_functions_0|redist10|delay_signals[1][28]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[0][28]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[0][28] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[0][28] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_36~0 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist10|delay_signals[0][28]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_36~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_36~0 .extended_lut = "off";
defparam \fp_functions_0|Mux_36~0 .lut_mask = 64'h0002000200020002;
defparam \fp_functions_0|Mux_36~0 .shared_arith = "off";

dffeas \fp_functions_0|redist10|delay_signals[0][29] (
	.clk(clk),
	.d(\fp_functions_0|redist10|delay_signals[1][29]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[0][29]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[0][29] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[0][29] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_35~0 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist10|delay_signals[0][29]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_35~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_35~0 .extended_lut = "off";
defparam \fp_functions_0|Mux_35~0 .lut_mask = 64'h0002000200020002;
defparam \fp_functions_0|Mux_35~0 .shared_arith = "off";

dffeas \fp_functions_0|redist10|delay_signals[0][30] (
	.clk(clk),
	.d(\fp_functions_0|redist10|delay_signals[1][30]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[0][30]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[0][30] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[0][30] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_34~0 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist10|delay_signals[0][30]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_34~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_34~0 .extended_lut = "off";
defparam \fp_functions_0|Mux_34~0 .lut_mask = 64'h0002000200020002;
defparam \fp_functions_0|Mux_34~0 .shared_arith = "off";

dffeas \fp_functions_0|redist10|delay_signals[0][31] (
	.clk(clk),
	.d(\fp_functions_0|redist10|delay_signals[1][31]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[0][31]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[0][31] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[0][31] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_33~0 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist10|delay_signals[0][31]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_33~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_33~0 .extended_lut = "off";
defparam \fp_functions_0|Mux_33~0 .lut_mask = 64'h0002000200020002;
defparam \fp_functions_0|Mux_33~0 .shared_arith = "off";

dffeas \fp_functions_0|redist10|delay_signals[0][32] (
	.clk(clk),
	.d(\fp_functions_0|redist10|delay_signals[1][32]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[0][32]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[0][32] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[0][32] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_32~0 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist10|delay_signals[0][32]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_32~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_32~0 .extended_lut = "off";
defparam \fp_functions_0|Mux_32~0 .lut_mask = 64'h0002000200020002;
defparam \fp_functions_0|Mux_32~0 .shared_arith = "off";

dffeas \fp_functions_0|redist10|delay_signals[0][33] (
	.clk(clk),
	.d(\fp_functions_0|redist10|delay_signals[1][33]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[0][33]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[0][33] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[0][33] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_31~0 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist10|delay_signals[0][33]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_31~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_31~0 .extended_lut = "off";
defparam \fp_functions_0|Mux_31~0 .lut_mask = 64'h0002000200020002;
defparam \fp_functions_0|Mux_31~0 .shared_arith = "off";

dffeas \fp_functions_0|redist10|delay_signals[0][34] (
	.clk(clk),
	.d(\fp_functions_0|redist10|delay_signals[1][34]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[0][34]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[0][34] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[0][34] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_30~0 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist10|delay_signals[0][34]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_30~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_30~0 .extended_lut = "off";
defparam \fp_functions_0|Mux_30~0 .lut_mask = 64'h0002000200020002;
defparam \fp_functions_0|Mux_30~0 .shared_arith = "off";

dffeas \fp_functions_0|redist10|delay_signals[0][35] (
	.clk(clk),
	.d(\fp_functions_0|redist10|delay_signals[1][35]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[0][35]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[0][35] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[0][35] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_29~0 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist10|delay_signals[0][35]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_29~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_29~0 .extended_lut = "off";
defparam \fp_functions_0|Mux_29~0 .lut_mask = 64'h0002000200020002;
defparam \fp_functions_0|Mux_29~0 .shared_arith = "off";

dffeas \fp_functions_0|redist10|delay_signals[0][36] (
	.clk(clk),
	.d(\fp_functions_0|redist10|delay_signals[1][36]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[0][36]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[0][36] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[0][36] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_28~0 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist10|delay_signals[0][36]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_28~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_28~0 .extended_lut = "off";
defparam \fp_functions_0|Mux_28~0 .lut_mask = 64'h0002000200020002;
defparam \fp_functions_0|Mux_28~0 .shared_arith = "off";

dffeas \fp_functions_0|redist10|delay_signals[0][37] (
	.clk(clk),
	.d(\fp_functions_0|redist10|delay_signals[1][37]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[0][37]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[0][37] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[0][37] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_27~0 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist10|delay_signals[0][37]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_27~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_27~0 .extended_lut = "off";
defparam \fp_functions_0|Mux_27~0 .lut_mask = 64'h0002000200020002;
defparam \fp_functions_0|Mux_27~0 .shared_arith = "off";

dffeas \fp_functions_0|redist10|delay_signals[0][38] (
	.clk(clk),
	.d(\fp_functions_0|redist10|delay_signals[1][38]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[0][38]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[0][38] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[0][38] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_26~0 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist10|delay_signals[0][38]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_26~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_26~0 .extended_lut = "off";
defparam \fp_functions_0|Mux_26~0 .lut_mask = 64'h0002000200020002;
defparam \fp_functions_0|Mux_26~0 .shared_arith = "off";

dffeas \fp_functions_0|redist10|delay_signals[0][39] (
	.clk(clk),
	.d(\fp_functions_0|redist10|delay_signals[1][39]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[0][39]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[0][39] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[0][39] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_25~0 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist10|delay_signals[0][39]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_25~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_25~0 .extended_lut = "off";
defparam \fp_functions_0|Mux_25~0 .lut_mask = 64'h0002000200020002;
defparam \fp_functions_0|Mux_25~0 .shared_arith = "off";

dffeas \fp_functions_0|redist10|delay_signals[0][40] (
	.clk(clk),
	.d(\fp_functions_0|redist10|delay_signals[1][40]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[0][40]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[0][40] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[0][40] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_24~0 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist10|delay_signals[0][40]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_24~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_24~0 .extended_lut = "off";
defparam \fp_functions_0|Mux_24~0 .lut_mask = 64'h0002000200020002;
defparam \fp_functions_0|Mux_24~0 .shared_arith = "off";

dffeas \fp_functions_0|redist10|delay_signals[0][41] (
	.clk(clk),
	.d(\fp_functions_0|redist10|delay_signals[1][41]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[0][41]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[0][41] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[0][41] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_23~0 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist10|delay_signals[0][41]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_23~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_23~0 .extended_lut = "off";
defparam \fp_functions_0|Mux_23~0 .lut_mask = 64'h0002000200020002;
defparam \fp_functions_0|Mux_23~0 .shared_arith = "off";

dffeas \fp_functions_0|redist10|delay_signals[0][42] (
	.clk(clk),
	.d(\fp_functions_0|redist10|delay_signals[1][42]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[0][42]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[0][42] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[0][42] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_22~0 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist10|delay_signals[0][42]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_22~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_22~0 .extended_lut = "off";
defparam \fp_functions_0|Mux_22~0 .lut_mask = 64'h0002000200020002;
defparam \fp_functions_0|Mux_22~0 .shared_arith = "off";

dffeas \fp_functions_0|redist10|delay_signals[0][43] (
	.clk(clk),
	.d(\fp_functions_0|redist10|delay_signals[1][43]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[0][43]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[0][43] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[0][43] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_21~0 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist10|delay_signals[0][43]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_21~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_21~0 .extended_lut = "off";
defparam \fp_functions_0|Mux_21~0 .lut_mask = 64'h0002000200020002;
defparam \fp_functions_0|Mux_21~0 .shared_arith = "off";

dffeas \fp_functions_0|redist10|delay_signals[0][44] (
	.clk(clk),
	.d(\fp_functions_0|redist10|delay_signals[1][44]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[0][44]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[0][44] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[0][44] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_20~0 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist10|delay_signals[0][44]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_20~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_20~0 .extended_lut = "off";
defparam \fp_functions_0|Mux_20~0 .lut_mask = 64'h0002000200020002;
defparam \fp_functions_0|Mux_20~0 .shared_arith = "off";

dffeas \fp_functions_0|redist10|delay_signals[0][45] (
	.clk(clk),
	.d(\fp_functions_0|redist10|delay_signals[1][45]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[0][45]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[0][45] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[0][45] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_19~0 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist10|delay_signals[0][45]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_19~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_19~0 .extended_lut = "off";
defparam \fp_functions_0|Mux_19~0 .lut_mask = 64'h0002000200020002;
defparam \fp_functions_0|Mux_19~0 .shared_arith = "off";

dffeas \fp_functions_0|redist10|delay_signals[0][46] (
	.clk(clk),
	.d(\fp_functions_0|redist10|delay_signals[1][46]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[0][46]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[0][46] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[0][46] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_18~0 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist10|delay_signals[0][46]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_18~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_18~0 .extended_lut = "off";
defparam \fp_functions_0|Mux_18~0 .lut_mask = 64'h0002000200020002;
defparam \fp_functions_0|Mux_18~0 .shared_arith = "off";

dffeas \fp_functions_0|redist10|delay_signals[0][47] (
	.clk(clk),
	.d(\fp_functions_0|redist10|delay_signals[1][47]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[0][47]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[0][47] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[0][47] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_17~0 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist10|delay_signals[0][47]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_17~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_17~0 .extended_lut = "off";
defparam \fp_functions_0|Mux_17~0 .lut_mask = 64'h0002000200020002;
defparam \fp_functions_0|Mux_17~0 .shared_arith = "off";

dffeas \fp_functions_0|redist10|delay_signals[0][48] (
	.clk(clk),
	.d(\fp_functions_0|redist10|delay_signals[1][48]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[0][48]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[0][48] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[0][48] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_16~0 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist10|delay_signals[0][48]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_16~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_16~0 .extended_lut = "off";
defparam \fp_functions_0|Mux_16~0 .lut_mask = 64'h0002000200020002;
defparam \fp_functions_0|Mux_16~0 .shared_arith = "off";

dffeas \fp_functions_0|redist10|delay_signals[0][49] (
	.clk(clk),
	.d(\fp_functions_0|redist10|delay_signals[1][49]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[0][49]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[0][49] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[0][49] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_15~0 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist10|delay_signals[0][49]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_15~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_15~0 .extended_lut = "off";
defparam \fp_functions_0|Mux_15~0 .lut_mask = 64'h0002000200020002;
defparam \fp_functions_0|Mux_15~0 .shared_arith = "off";

dffeas \fp_functions_0|redist10|delay_signals[0][50] (
	.clk(clk),
	.d(\fp_functions_0|redist10|delay_signals[1][50]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[0][50]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[0][50] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[0][50] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_14~0 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist10|delay_signals[0][50]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_14~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_14~0 .extended_lut = "off";
defparam \fp_functions_0|Mux_14~0 .lut_mask = 64'h0002000200020002;
defparam \fp_functions_0|Mux_14~0 .shared_arith = "off";

dffeas \fp_functions_0|redist10|delay_signals[0][51] (
	.clk(clk),
	.d(\fp_functions_0|redist10|delay_signals[1][51]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[0][51]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[0][51] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[0][51] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_13~0 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist10|delay_signals[0][51]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_13~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_13~0 .extended_lut = "off";
defparam \fp_functions_0|Mux_13~0 .lut_mask = 64'h0002000200020002;
defparam \fp_functions_0|Mux_13~0 .shared_arith = "off";

dffeas \fp_functions_0|redist8|delay_signals[0][0] (
	.clk(clk),
	.d(\fp_functions_0|redist9|delay_signals[0][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist8|delay_signals[0][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist8|delay_signals[0][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist8|delay_signals[0][0] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_12~0 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist8|delay_signals[0][0]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_12~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_12~0 .extended_lut = "off";
defparam \fp_functions_0|Mux_12~0 .lut_mask = 64'h00A700A700A700A7;
defparam \fp_functions_0|Mux_12~0 .shared_arith = "off";

dffeas \fp_functions_0|redist8|delay_signals[0][1] (
	.clk(clk),
	.d(\fp_functions_0|redist9|delay_signals[0][1]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist8|delay_signals[0][1]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist8|delay_signals[0][1] .is_wysiwyg = "true";
defparam \fp_functions_0|redist8|delay_signals[0][1] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_12~1 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist8|delay_signals[0][1]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_12~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_12~1 .extended_lut = "off";
defparam \fp_functions_0|Mux_12~1 .lut_mask = 64'h00A700A700A700A7;
defparam \fp_functions_0|Mux_12~1 .shared_arith = "off";

dffeas \fp_functions_0|redist8|delay_signals[0][2] (
	.clk(clk),
	.d(\fp_functions_0|redist9|delay_signals[0][2]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist8|delay_signals[0][2]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist8|delay_signals[0][2] .is_wysiwyg = "true";
defparam \fp_functions_0|redist8|delay_signals[0][2] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_12~2 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist8|delay_signals[0][2]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_12~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_12~2 .extended_lut = "off";
defparam \fp_functions_0|Mux_12~2 .lut_mask = 64'h00A700A700A700A7;
defparam \fp_functions_0|Mux_12~2 .shared_arith = "off";

dffeas \fp_functions_0|redist8|delay_signals[0][3] (
	.clk(clk),
	.d(\fp_functions_0|redist9|delay_signals[0][3]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist8|delay_signals[0][3]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist8|delay_signals[0][3] .is_wysiwyg = "true";
defparam \fp_functions_0|redist8|delay_signals[0][3] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_12~3 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist8|delay_signals[0][3]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_12~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_12~3 .extended_lut = "off";
defparam \fp_functions_0|Mux_12~3 .lut_mask = 64'h00A700A700A700A7;
defparam \fp_functions_0|Mux_12~3 .shared_arith = "off";

dffeas \fp_functions_0|redist8|delay_signals[0][4] (
	.clk(clk),
	.d(\fp_functions_0|redist9|delay_signals[0][4]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist8|delay_signals[0][4]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist8|delay_signals[0][4] .is_wysiwyg = "true";
defparam \fp_functions_0|redist8|delay_signals[0][4] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_12~4 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist8|delay_signals[0][4]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_12~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_12~4 .extended_lut = "off";
defparam \fp_functions_0|Mux_12~4 .lut_mask = 64'h00A700A700A700A7;
defparam \fp_functions_0|Mux_12~4 .shared_arith = "off";

dffeas \fp_functions_0|redist8|delay_signals[0][5] (
	.clk(clk),
	.d(\fp_functions_0|redist9|delay_signals[0][5]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist8|delay_signals[0][5]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist8|delay_signals[0][5] .is_wysiwyg = "true";
defparam \fp_functions_0|redist8|delay_signals[0][5] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_12~5 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist8|delay_signals[0][5]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_12~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_12~5 .extended_lut = "off";
defparam \fp_functions_0|Mux_12~5 .lut_mask = 64'h00A700A700A700A7;
defparam \fp_functions_0|Mux_12~5 .shared_arith = "off";

dffeas \fp_functions_0|redist8|delay_signals[0][6] (
	.clk(clk),
	.d(\fp_functions_0|redist9|delay_signals[0][6]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist8|delay_signals[0][6]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist8|delay_signals[0][6] .is_wysiwyg = "true";
defparam \fp_functions_0|redist8|delay_signals[0][6] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_12~6 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist8|delay_signals[0][6]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_12~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_12~6 .extended_lut = "off";
defparam \fp_functions_0|Mux_12~6 .lut_mask = 64'h00A700A700A700A7;
defparam \fp_functions_0|Mux_12~6 .shared_arith = "off";

dffeas \fp_functions_0|redist8|delay_signals[0][7] (
	.clk(clk),
	.d(\fp_functions_0|redist9|delay_signals[0][7]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist8|delay_signals[0][7]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist8|delay_signals[0][7] .is_wysiwyg = "true";
defparam \fp_functions_0|redist8|delay_signals[0][7] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_12~7 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist8|delay_signals[0][7]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_12~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_12~7 .extended_lut = "off";
defparam \fp_functions_0|Mux_12~7 .lut_mask = 64'h00A700A700A700A7;
defparam \fp_functions_0|Mux_12~7 .shared_arith = "off";

dffeas \fp_functions_0|redist8|delay_signals[0][8] (
	.clk(clk),
	.d(\fp_functions_0|redist9|delay_signals[0][8]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist8|delay_signals[0][8]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist8|delay_signals[0][8] .is_wysiwyg = "true";
defparam \fp_functions_0|redist8|delay_signals[0][8] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_12~8 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist8|delay_signals[0][8]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_12~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_12~8 .extended_lut = "off";
defparam \fp_functions_0|Mux_12~8 .lut_mask = 64'h00A700A700A700A7;
defparam \fp_functions_0|Mux_12~8 .shared_arith = "off";

dffeas \fp_functions_0|redist8|delay_signals[0][9] (
	.clk(clk),
	.d(\fp_functions_0|redist9|delay_signals[0][9]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist8|delay_signals[0][9]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist8|delay_signals[0][9] .is_wysiwyg = "true";
defparam \fp_functions_0|redist8|delay_signals[0][9] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_12~9 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist8|delay_signals[0][9]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_12~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_12~9 .extended_lut = "off";
defparam \fp_functions_0|Mux_12~9 .lut_mask = 64'h00A700A700A700A7;
defparam \fp_functions_0|Mux_12~9 .shared_arith = "off";

dffeas \fp_functions_0|redist8|delay_signals[0][10] (
	.clk(clk),
	.d(\fp_functions_0|redist9|delay_signals[0][10]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist8|delay_signals[0][10]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist8|delay_signals[0][10] .is_wysiwyg = "true";
defparam \fp_functions_0|redist8|delay_signals[0][10] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|Mux_12~10 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist8|delay_signals[0][10]~q ),
	.datac(!\fp_functions_0|i6400~combout ),
	.datad(!\fp_functions_0|i6475~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|Mux_12~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|Mux_12~10 .extended_lut = "off";
defparam \fp_functions_0|Mux_12~10 .lut_mask = 64'h00A700A700A700A7;
defparam \fp_functions_0|Mux_12~10 .shared_arith = "off";

dffeas \fp_functions_0|redist14|delay_signals[0][0] (
	.clk(clk),
	.d(\fp_functions_0|redist14|delay_signals[1][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist14|delay_signals[0][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist14|delay_signals[0][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist14|delay_signals[0][0] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|i1071 (
	.dataa(!\fp_functions_0|excRNaN_uid89_fpMulTest_delay|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist14|delay_signals[0][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|i1071~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|i1071 .extended_lut = "off";
defparam \fp_functions_0|i1071 .lut_mask = 64'h2222222222222222;
defparam \fp_functions_0|i1071 .shared_arith = "off";

dffeas \fp_functions_0|redist10|delay_signals[1][0] (
	.clk(clk),
	.d(\fp_functions_0|add_6~1_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[1][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[1][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[1][0] .power_up = "low";

dffeas \fp_functions_0|redist18|delay_signals[0][0] (
	.clk(clk),
	.d(\fp_functions_0|redist18|delay_signals[1][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist18|delay_signals[0][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist18|delay_signals[0][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist18|delay_signals[0][0] .power_up = "low";

dffeas \fp_functions_0|redist17|delay_signals[0][0] (
	.clk(clk),
	.d(\fp_functions_0|redist17|delay_signals[1][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist17|delay_signals[0][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist17|delay_signals[0][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist17|delay_signals[0][0] .power_up = "low";

dffeas \fp_functions_0|redist20|delay_signals[0][0] (
	.clk(clk),
	.d(\fp_functions_0|redist20|delay_signals[1][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist20|delay_signals[0][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist20|delay_signals[0][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist20|delay_signals[0][0] .power_up = "low";

dffeas \fp_functions_0|redist21|delay_signals[0][0] (
	.clk(clk),
	.d(\fp_functions_0|redist21|delay_signals[1][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist21|delay_signals[0][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist21|delay_signals[0][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist21|delay_signals[0][0] .power_up = "low";

dffeas \fp_functions_0|redist16|delay_signals[0][0] (
	.clk(clk),
	.d(\fp_functions_0|redist16|delay_signals[1][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist16|delay_signals[0][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist16|delay_signals[0][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist16|delay_signals[0][0] .power_up = "low";

dffeas \fp_functions_0|redist19|delay_signals[0][0] (
	.clk(clk),
	.d(\fp_functions_0|redist19|delay_signals[1][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist19|delay_signals[0][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist19|delay_signals[0][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist19|delay_signals[0][0] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|i933~0 (
	.dataa(!\fp_functions_0|redist18|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist17|delay_signals[0][0]~q ),
	.datac(!\fp_functions_0|redist20|delay_signals[0][0]~q ),
	.datad(!\fp_functions_0|redist21|delay_signals[0][0]~q ),
	.datae(!\fp_functions_0|redist16|delay_signals[0][0]~q ),
	.dataf(!\fp_functions_0|redist19|delay_signals[0][0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|i933~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|i933~0 .extended_lut = "off";
defparam \fp_functions_0|i933~0 .lut_mask = 64'h3F3F0F3F37370537;
defparam \fp_functions_0|i933~0 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|i6384 (
	.dataa(!\fp_functions_0|redist18|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist17|delay_signals[0][0]~q ),
	.datac(!\fp_functions_0|redist20|delay_signals[0][0]~q ),
	.datad(!\fp_functions_0|redist21|delay_signals[0][0]~q ),
	.datae(!\fp_functions_0|add_7~1_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|i6384~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|i6384 .extended_lut = "off";
defparam \fp_functions_0|i6384 .lut_mask = 64'h8000000080000000;
defparam \fp_functions_0|i6384 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|i6387~0 (
	.dataa(!\fp_functions_0|redist18|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist17|delay_signals[0][0]~q ),
	.datac(!\fp_functions_0|redist20|delay_signals[0][0]~q ),
	.datad(!\fp_functions_0|redist19|delay_signals[0][0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|i6387~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|i6387~0 .extended_lut = "off";
defparam \fp_functions_0|i6387~0 .lut_mask = 64'h0008000800080008;
defparam \fp_functions_0|i6387~0 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|i6390~0 (
	.dataa(!\fp_functions_0|redist17|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist20|delay_signals[0][0]~q ),
	.datac(!\fp_functions_0|redist21|delay_signals[0][0]~q ),
	.datad(!\fp_functions_0|redist16|delay_signals[0][0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|i6390~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|i6390~0 .extended_lut = "off";
defparam \fp_functions_0|i6390~0 .lut_mask = 64'h0040004000400040;
defparam \fp_functions_0|i6390~0 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|i6393~0 (
	.dataa(!\fp_functions_0|redist17|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist20|delay_signals[0][0]~q ),
	.datac(!\fp_functions_0|redist16|delay_signals[0][0]~q ),
	.datad(!\fp_functions_0|redist19|delay_signals[0][0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|i6393~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|i6393~0 .extended_lut = "off";
defparam \fp_functions_0|i6393~0 .lut_mask = 64'h0001000100010001;
defparam \fp_functions_0|i6393~0 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|i6459 (
	.dataa(!\fp_functions_0|redist18|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist17|delay_signals[0][0]~q ),
	.datac(!\fp_functions_0|redist20|delay_signals[0][0]~q ),
	.datad(!\fp_functions_0|redist21|delay_signals[0][0]~q ),
	.datae(!\fp_functions_0|add_8~1_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|i6459~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|i6459 .extended_lut = "off";
defparam \fp_functions_0|i6459 .lut_mask = 64'h8000000080000000;
defparam \fp_functions_0|i6459 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|i6462~0 (
	.dataa(!\fp_functions_0|redist18|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist20|delay_signals[0][0]~q ),
	.datac(!\fp_functions_0|redist21|delay_signals[0][0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|i6462~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|i6462~0 .extended_lut = "off";
defparam \fp_functions_0|i6462~0 .lut_mask = 64'h4040404040404040;
defparam \fp_functions_0|i6462~0 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|i6465~0 (
	.dataa(!\fp_functions_0|redist18|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist17|delay_signals[0][0]~q ),
	.datac(!\fp_functions_0|redist21|delay_signals[0][0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|i6465~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|i6465~0 .extended_lut = "off";
defparam \fp_functions_0|i6465~0 .lut_mask = 64'h0808080808080808;
defparam \fp_functions_0|i6465~0 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|i6468 (
	.dataa(!\fp_functions_0|redist18|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist21|delay_signals[0][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|i6468~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|i6468 .extended_lut = "off";
defparam \fp_functions_0|i6468 .lut_mask = 64'h1111111111111111;
defparam \fp_functions_0|i6468 .shared_arith = "off";

dffeas \fp_functions_0|redist10|delay_signals[1][1] (
	.clk(clk),
	.d(\fp_functions_0|add_6~5_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[1][1]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[1][1] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[1][1] .power_up = "low";

dffeas \fp_functions_0|redist10|delay_signals[1][2] (
	.clk(clk),
	.d(\fp_functions_0|add_6~9_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[1][2]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[1][2] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[1][2] .power_up = "low";

dffeas \fp_functions_0|redist10|delay_signals[1][3] (
	.clk(clk),
	.d(\fp_functions_0|add_6~13_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[1][3]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[1][3] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[1][3] .power_up = "low";

dffeas \fp_functions_0|redist10|delay_signals[1][4] (
	.clk(clk),
	.d(\fp_functions_0|add_6~17_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[1][4]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[1][4] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[1][4] .power_up = "low";

dffeas \fp_functions_0|redist10|delay_signals[1][5] (
	.clk(clk),
	.d(\fp_functions_0|add_6~21_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[1][5]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[1][5] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[1][5] .power_up = "low";

dffeas \fp_functions_0|redist10|delay_signals[1][6] (
	.clk(clk),
	.d(\fp_functions_0|add_6~25_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[1][6]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[1][6] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[1][6] .power_up = "low";

dffeas \fp_functions_0|redist10|delay_signals[1][7] (
	.clk(clk),
	.d(\fp_functions_0|add_6~29_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[1][7]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[1][7] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[1][7] .power_up = "low";

dffeas \fp_functions_0|redist10|delay_signals[1][8] (
	.clk(clk),
	.d(\fp_functions_0|add_6~33_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[1][8]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[1][8] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[1][8] .power_up = "low";

dffeas \fp_functions_0|redist10|delay_signals[1][9] (
	.clk(clk),
	.d(\fp_functions_0|add_6~37_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[1][9]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[1][9] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[1][9] .power_up = "low";

dffeas \fp_functions_0|redist10|delay_signals[1][10] (
	.clk(clk),
	.d(\fp_functions_0|add_6~41_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[1][10]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[1][10] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[1][10] .power_up = "low";

dffeas \fp_functions_0|redist10|delay_signals[1][11] (
	.clk(clk),
	.d(\fp_functions_0|add_6~45_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[1][11]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[1][11] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[1][11] .power_up = "low";

dffeas \fp_functions_0|redist10|delay_signals[1][12] (
	.clk(clk),
	.d(\fp_functions_0|add_6~49_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[1][12]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[1][12] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[1][12] .power_up = "low";

dffeas \fp_functions_0|redist10|delay_signals[1][13] (
	.clk(clk),
	.d(\fp_functions_0|add_6~53_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[1][13]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[1][13] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[1][13] .power_up = "low";

dffeas \fp_functions_0|redist10|delay_signals[1][14] (
	.clk(clk),
	.d(\fp_functions_0|add_6~57_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[1][14]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[1][14] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[1][14] .power_up = "low";

dffeas \fp_functions_0|redist10|delay_signals[1][15] (
	.clk(clk),
	.d(\fp_functions_0|add_6~61_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[1][15]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[1][15] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[1][15] .power_up = "low";

dffeas \fp_functions_0|redist10|delay_signals[1][16] (
	.clk(clk),
	.d(\fp_functions_0|add_6~65_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[1][16]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[1][16] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[1][16] .power_up = "low";

dffeas \fp_functions_0|redist10|delay_signals[1][17] (
	.clk(clk),
	.d(\fp_functions_0|add_6~69_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[1][17]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[1][17] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[1][17] .power_up = "low";

dffeas \fp_functions_0|redist10|delay_signals[1][18] (
	.clk(clk),
	.d(\fp_functions_0|add_6~73_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[1][18]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[1][18] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[1][18] .power_up = "low";

dffeas \fp_functions_0|redist10|delay_signals[1][19] (
	.clk(clk),
	.d(\fp_functions_0|add_6~77_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[1][19]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[1][19] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[1][19] .power_up = "low";

dffeas \fp_functions_0|redist10|delay_signals[1][20] (
	.clk(clk),
	.d(\fp_functions_0|add_6~81_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[1][20]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[1][20] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[1][20] .power_up = "low";

dffeas \fp_functions_0|redist10|delay_signals[1][21] (
	.clk(clk),
	.d(\fp_functions_0|add_6~85_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[1][21]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[1][21] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[1][21] .power_up = "low";

dffeas \fp_functions_0|redist10|delay_signals[1][22] (
	.clk(clk),
	.d(\fp_functions_0|add_6~89_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[1][22]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[1][22] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[1][22] .power_up = "low";

dffeas \fp_functions_0|redist10|delay_signals[1][23] (
	.clk(clk),
	.d(\fp_functions_0|add_6~93_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[1][23]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[1][23] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[1][23] .power_up = "low";

dffeas \fp_functions_0|redist10|delay_signals[1][24] (
	.clk(clk),
	.d(\fp_functions_0|add_6~97_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[1][24]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[1][24] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[1][24] .power_up = "low";

dffeas \fp_functions_0|redist10|delay_signals[1][25] (
	.clk(clk),
	.d(\fp_functions_0|add_6~101_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[1][25]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[1][25] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[1][25] .power_up = "low";

dffeas \fp_functions_0|redist10|delay_signals[1][26] (
	.clk(clk),
	.d(\fp_functions_0|add_6~105_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[1][26]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[1][26] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[1][26] .power_up = "low";

dffeas \fp_functions_0|redist10|delay_signals[1][27] (
	.clk(clk),
	.d(\fp_functions_0|add_6~109_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[1][27]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[1][27] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[1][27] .power_up = "low";

dffeas \fp_functions_0|redist10|delay_signals[1][28] (
	.clk(clk),
	.d(\fp_functions_0|add_6~113_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[1][28]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[1][28] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[1][28] .power_up = "low";

dffeas \fp_functions_0|redist10|delay_signals[1][29] (
	.clk(clk),
	.d(\fp_functions_0|add_6~117_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[1][29]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[1][29] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[1][29] .power_up = "low";

dffeas \fp_functions_0|redist10|delay_signals[1][30] (
	.clk(clk),
	.d(\fp_functions_0|add_6~121_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[1][30]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[1][30] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[1][30] .power_up = "low";

dffeas \fp_functions_0|redist10|delay_signals[1][31] (
	.clk(clk),
	.d(\fp_functions_0|add_6~125_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[1][31]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[1][31] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[1][31] .power_up = "low";

dffeas \fp_functions_0|redist10|delay_signals[1][32] (
	.clk(clk),
	.d(\fp_functions_0|add_6~129_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[1][32]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[1][32] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[1][32] .power_up = "low";

dffeas \fp_functions_0|redist10|delay_signals[1][33] (
	.clk(clk),
	.d(\fp_functions_0|add_6~133_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[1][33]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[1][33] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[1][33] .power_up = "low";

dffeas \fp_functions_0|redist10|delay_signals[1][34] (
	.clk(clk),
	.d(\fp_functions_0|add_6~137_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[1][34]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[1][34] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[1][34] .power_up = "low";

dffeas \fp_functions_0|redist10|delay_signals[1][35] (
	.clk(clk),
	.d(\fp_functions_0|add_6~141_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[1][35]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[1][35] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[1][35] .power_up = "low";

dffeas \fp_functions_0|redist10|delay_signals[1][36] (
	.clk(clk),
	.d(\fp_functions_0|add_6~145_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[1][36]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[1][36] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[1][36] .power_up = "low";

dffeas \fp_functions_0|redist10|delay_signals[1][37] (
	.clk(clk),
	.d(\fp_functions_0|add_6~149_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[1][37]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[1][37] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[1][37] .power_up = "low";

dffeas \fp_functions_0|redist10|delay_signals[1][38] (
	.clk(clk),
	.d(\fp_functions_0|add_6~153_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[1][38]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[1][38] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[1][38] .power_up = "low";

dffeas \fp_functions_0|redist10|delay_signals[1][39] (
	.clk(clk),
	.d(\fp_functions_0|add_6~157_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[1][39]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[1][39] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[1][39] .power_up = "low";

dffeas \fp_functions_0|redist10|delay_signals[1][40] (
	.clk(clk),
	.d(\fp_functions_0|add_6~161_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[1][40]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[1][40] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[1][40] .power_up = "low";

dffeas \fp_functions_0|redist10|delay_signals[1][41] (
	.clk(clk),
	.d(\fp_functions_0|add_6~165_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[1][41]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[1][41] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[1][41] .power_up = "low";

dffeas \fp_functions_0|redist10|delay_signals[1][42] (
	.clk(clk),
	.d(\fp_functions_0|add_6~169_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[1][42]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[1][42] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[1][42] .power_up = "low";

dffeas \fp_functions_0|redist10|delay_signals[1][43] (
	.clk(clk),
	.d(\fp_functions_0|add_6~173_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[1][43]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[1][43] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[1][43] .power_up = "low";

dffeas \fp_functions_0|redist10|delay_signals[1][44] (
	.clk(clk),
	.d(\fp_functions_0|add_6~177_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[1][44]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[1][44] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[1][44] .power_up = "low";

dffeas \fp_functions_0|redist10|delay_signals[1][45] (
	.clk(clk),
	.d(\fp_functions_0|add_6~181_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[1][45]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[1][45] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[1][45] .power_up = "low";

dffeas \fp_functions_0|redist10|delay_signals[1][46] (
	.clk(clk),
	.d(\fp_functions_0|add_6~185_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[1][46]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[1][46] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[1][46] .power_up = "low";

dffeas \fp_functions_0|redist10|delay_signals[1][47] (
	.clk(clk),
	.d(\fp_functions_0|add_6~189_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[1][47]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[1][47] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[1][47] .power_up = "low";

dffeas \fp_functions_0|redist10|delay_signals[1][48] (
	.clk(clk),
	.d(\fp_functions_0|add_6~193_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[1][48]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[1][48] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[1][48] .power_up = "low";

dffeas \fp_functions_0|redist10|delay_signals[1][49] (
	.clk(clk),
	.d(\fp_functions_0|add_6~197_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[1][49]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[1][49] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[1][49] .power_up = "low";

dffeas \fp_functions_0|redist10|delay_signals[1][50] (
	.clk(clk),
	.d(\fp_functions_0|add_6~201_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[1][50]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[1][50] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[1][50] .power_up = "low";

dffeas \fp_functions_0|redist10|delay_signals[1][51] (
	.clk(clk),
	.d(\fp_functions_0|add_6~205_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist10|delay_signals[1][51]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist10|delay_signals[1][51] .is_wysiwyg = "true";
defparam \fp_functions_0|redist10|delay_signals[1][51] .power_up = "low";

dffeas \fp_functions_0|redist9|delay_signals[0][0] (
	.clk(clk),
	.d(\fp_functions_0|add_6~209_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist9|delay_signals[0][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist9|delay_signals[0][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist9|delay_signals[0][0] .power_up = "low";

dffeas \fp_functions_0|redist9|delay_signals[0][1] (
	.clk(clk),
	.d(\fp_functions_0|add_6~213_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist9|delay_signals[0][1]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist9|delay_signals[0][1] .is_wysiwyg = "true";
defparam \fp_functions_0|redist9|delay_signals[0][1] .power_up = "low";

dffeas \fp_functions_0|redist9|delay_signals[0][2] (
	.clk(clk),
	.d(\fp_functions_0|add_6~217_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist9|delay_signals[0][2]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist9|delay_signals[0][2] .is_wysiwyg = "true";
defparam \fp_functions_0|redist9|delay_signals[0][2] .power_up = "low";

dffeas \fp_functions_0|redist9|delay_signals[0][3] (
	.clk(clk),
	.d(\fp_functions_0|add_6~221_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist9|delay_signals[0][3]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist9|delay_signals[0][3] .is_wysiwyg = "true";
defparam \fp_functions_0|redist9|delay_signals[0][3] .power_up = "low";

dffeas \fp_functions_0|redist9|delay_signals[0][4] (
	.clk(clk),
	.d(\fp_functions_0|add_6~225_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist9|delay_signals[0][4]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist9|delay_signals[0][4] .is_wysiwyg = "true";
defparam \fp_functions_0|redist9|delay_signals[0][4] .power_up = "low";

dffeas \fp_functions_0|redist9|delay_signals[0][5] (
	.clk(clk),
	.d(\fp_functions_0|add_6~229_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist9|delay_signals[0][5]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist9|delay_signals[0][5] .is_wysiwyg = "true";
defparam \fp_functions_0|redist9|delay_signals[0][5] .power_up = "low";

dffeas \fp_functions_0|redist9|delay_signals[0][6] (
	.clk(clk),
	.d(\fp_functions_0|add_6~233_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist9|delay_signals[0][6]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist9|delay_signals[0][6] .is_wysiwyg = "true";
defparam \fp_functions_0|redist9|delay_signals[0][6] .power_up = "low";

dffeas \fp_functions_0|redist9|delay_signals[0][7] (
	.clk(clk),
	.d(\fp_functions_0|add_6~237_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist9|delay_signals[0][7]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist9|delay_signals[0][7] .is_wysiwyg = "true";
defparam \fp_functions_0|redist9|delay_signals[0][7] .power_up = "low";

dffeas \fp_functions_0|redist9|delay_signals[0][8] (
	.clk(clk),
	.d(\fp_functions_0|add_6~241_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist9|delay_signals[0][8]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist9|delay_signals[0][8] .is_wysiwyg = "true";
defparam \fp_functions_0|redist9|delay_signals[0][8] .power_up = "low";

dffeas \fp_functions_0|redist9|delay_signals[0][9] (
	.clk(clk),
	.d(\fp_functions_0|add_6~245_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist9|delay_signals[0][9]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist9|delay_signals[0][9] .is_wysiwyg = "true";
defparam \fp_functions_0|redist9|delay_signals[0][9] .power_up = "low";

dffeas \fp_functions_0|redist9|delay_signals[0][10] (
	.clk(clk),
	.d(\fp_functions_0|add_6~249_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist9|delay_signals[0][10]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist9|delay_signals[0][10] .is_wysiwyg = "true";
defparam \fp_functions_0|redist9|delay_signals[0][10] .power_up = "low";

dffeas \fp_functions_0|redist14|delay_signals[1][0] (
	.clk(clk),
	.d(\fp_functions_0|redist14|delay_signals[2][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist14|delay_signals[1][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist14|delay_signals[1][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist14|delay_signals[1][0] .power_up = "low";

dffeas \fp_functions_0|redist18|delay_signals[1][0] (
	.clk(clk),
	.d(\fp_functions_0|redist18|delay_signals[2][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist18|delay_signals[1][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist18|delay_signals[1][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist18|delay_signals[1][0] .power_up = "low";

dffeas \fp_functions_0|redist17|delay_signals[1][0] (
	.clk(clk),
	.d(\fp_functions_0|redist17|delay_signals[2][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist17|delay_signals[1][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist17|delay_signals[1][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist17|delay_signals[1][0] .power_up = "low";

dffeas \fp_functions_0|redist20|delay_signals[1][0] (
	.clk(clk),
	.d(\fp_functions_0|redist20|delay_signals[2][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist20|delay_signals[1][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist20|delay_signals[1][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist20|delay_signals[1][0] .power_up = "low";

dffeas \fp_functions_0|redist21|delay_signals[1][0] (
	.clk(clk),
	.d(\fp_functions_0|redist21|delay_signals[2][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist21|delay_signals[1][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist21|delay_signals[1][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist21|delay_signals[1][0] .power_up = "low";

dffeas \fp_functions_0|redist16|delay_signals[1][0] (
	.clk(clk),
	.d(\fp_functions_0|redist16|delay_signals[2][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist16|delay_signals[1][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist16|delay_signals[1][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist16|delay_signals[1][0] .power_up = "low";

dffeas \fp_functions_0|redist19|delay_signals[1][0] (
	.clk(clk),
	.d(\fp_functions_0|redist19|delay_signals[2][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist19|delay_signals[1][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist19|delay_signals[1][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist19|delay_signals[1][0] .power_up = "low";

dffeas \fp_functions_0|redist9|delay_signals[0][14] (
	.clk(clk),
	.d(\fp_functions_0|add_6~257_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist9|delay_signals[0][14]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist9|delay_signals[0][14] .is_wysiwyg = "true";
defparam \fp_functions_0|redist9|delay_signals[0][14] .power_up = "low";

dffeas \fp_functions_0|redist14|delay_signals[2][0] (
	.clk(clk),
	.d(\fp_functions_0|redist14|delay_signals[3][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist14|delay_signals[2][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist14|delay_signals[2][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist14|delay_signals[2][0] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][1] (
	.clk(clk),
	.d(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[1]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][1]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][1] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][1] .power_up = "low";

dffeas \fp_functions_0|redist18|delay_signals[2][0] (
	.clk(clk),
	.d(\fp_functions_0|redist18|delay_signals[3][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist18|delay_signals[2][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist18|delay_signals[2][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist18|delay_signals[2][0] .power_up = "low";

dffeas \fp_functions_0|redist17|delay_signals[2][0] (
	.clk(clk),
	.d(\fp_functions_0|redist17|delay_signals[3][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist17|delay_signals[2][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist17|delay_signals[2][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist17|delay_signals[2][0] .power_up = "low";

dffeas \fp_functions_0|redist20|delay_signals[2][0] (
	.clk(clk),
	.d(\fp_functions_0|redist20|delay_signals[3][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist20|delay_signals[2][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist20|delay_signals[2][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist20|delay_signals[2][0] .power_up = "low";

dffeas \fp_functions_0|redist21|delay_signals[2][0] (
	.clk(clk),
	.d(\fp_functions_0|redist21|delay_signals[3][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist21|delay_signals[2][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist21|delay_signals[2][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist21|delay_signals[2][0] .power_up = "low";

dffeas \fp_functions_0|redist16|delay_signals[2][0] (
	.clk(clk),
	.d(\fp_functions_0|redist16|delay_signals[3][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist16|delay_signals[2][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist16|delay_signals[2][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist16|delay_signals[2][0] .power_up = "low";

dffeas \fp_functions_0|redist19|delay_signals[2][0] (
	.clk(clk),
	.d(\fp_functions_0|redist19|delay_signals[3][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist19|delay_signals[2][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist19|delay_signals[2][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist19|delay_signals[2][0] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][2] (
	.clk(clk),
	.d(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[2]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][2]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][2] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][2] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][3] (
	.clk(clk),
	.d(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[3]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][3]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][3] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][3] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][4] (
	.clk(clk),
	.d(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[4]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][4]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][4] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][4] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][5] (
	.clk(clk),
	.d(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[5]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][5]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][5] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][5] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][6] (
	.clk(clk),
	.d(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[6]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][6]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][6] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][6] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][7] (
	.clk(clk),
	.d(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[7]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][7]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][7] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][7] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][8] (
	.clk(clk),
	.d(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[8]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][8]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][8] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][8] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][9] (
	.clk(clk),
	.d(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[9]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][9]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][9] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][9] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][10] (
	.clk(clk),
	.d(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[10]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][10]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][10] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][10] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][11] (
	.clk(clk),
	.d(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[11]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][11]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][11] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][11] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][12] (
	.clk(clk),
	.d(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[12]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][12]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][12] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][12] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][13] (
	.clk(clk),
	.d(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[13]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][13]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][13] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][13] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][14] (
	.clk(clk),
	.d(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[14]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][14]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][14] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][14] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][15] (
	.clk(clk),
	.d(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[15]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][15]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][15] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][15] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][16] (
	.clk(clk),
	.d(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[16]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][16]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][16] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][16] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][17] (
	.clk(clk),
	.d(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[17]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][17]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][17] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][17] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][18] (
	.clk(clk),
	.d(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[18]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][18]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][18] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][18] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][19] (
	.clk(clk),
	.d(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[19]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][19]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][19] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][19] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][20] (
	.clk(clk),
	.d(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[20]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][20]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][20] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][20] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][21] (
	.clk(clk),
	.d(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[21]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][21]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][21] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][21] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][22] (
	.clk(clk),
	.d(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[22]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][22]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][22] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][22] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][23] (
	.clk(clk),
	.d(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[23]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][23]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][23] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][23] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][24] (
	.clk(clk),
	.d(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[24]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][24]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][24] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][24] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][25] (
	.clk(clk),
	.d(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[25]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][25]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][25] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][25] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][26] (
	.clk(clk),
	.d(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[26]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][26]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][26] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][26] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][27] (
	.clk(clk),
	.d(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[27]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][27]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][27] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][27] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][28] (
	.clk(clk),
	.d(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[28]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][28]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][28] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][28] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][29] (
	.clk(clk),
	.d(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[29]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][29]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][29] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][29] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][30] (
	.clk(clk),
	.d(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[30]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][30]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][30] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][30] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][31] (
	.clk(clk),
	.d(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[31]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][31]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][31] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][31] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][32] (
	.clk(clk),
	.d(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[32]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][32]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][32] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][32] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][33] (
	.clk(clk),
	.d(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[33]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][33]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][33] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][33] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][34] (
	.clk(clk),
	.d(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[34]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][34]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][34] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][34] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][35] (
	.clk(clk),
	.d(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[35]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][35]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][35] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][35] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][36] (
	.clk(clk),
	.d(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[36]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][36]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][36] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][36] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][37] (
	.clk(clk),
	.d(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[37]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][37]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][37] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][37] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][38] (
	.clk(clk),
	.d(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[38]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][38]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][38] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][38] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][39] (
	.clk(clk),
	.d(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[39]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][39]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][39] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][39] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][40] (
	.clk(clk),
	.d(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[40]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][40]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][40] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][40] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][41] (
	.clk(clk),
	.d(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[41]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][41]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][41] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][41] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][42] (
	.clk(clk),
	.d(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[42]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][42]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][42] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][42] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][43] (
	.clk(clk),
	.d(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[43]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][43]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][43] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][43] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][44] (
	.clk(clk),
	.d(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[44]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][44]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][44] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][44] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][45] (
	.clk(clk),
	.d(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[45]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][45]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][45] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][45] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][46] (
	.clk(clk),
	.d(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[46]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][46]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][46] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][46] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][47] (
	.clk(clk),
	.d(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[47]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][47]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][47] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][47] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][48] (
	.clk(clk),
	.d(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[48]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][48]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][48] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][48] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][49] (
	.clk(clk),
	.d(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[49]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][49]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][49] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][49] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][50] (
	.clk(clk),
	.d(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[50]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][50]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][50] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][50] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][51] (
	.clk(clk),
	.d(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[51]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][51]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][51] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][51] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][52] (
	.clk(clk),
	.d(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[52]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][52]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][52] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][52] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][53] (
	.clk(clk),
	.d(\fp_functions_0|redist11|delay_signals[0][53]~0_combout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][53]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][53] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][53] .power_up = "low";

dffeas \fp_functions_0|redist13|delay_signals[0][0] (
	.clk(clk),
	.d(\fp_functions_0|redist13|delay_signals[1][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist13|delay_signals[0][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist13|delay_signals[0][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist13|delay_signals[0][0] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][54] (
	.clk(clk),
	.d(\fp_functions_0|add_5~1_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][54]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][54] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][54] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][55] (
	.clk(clk),
	.d(\fp_functions_0|add_5~5_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][55]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][55] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][55] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][56] (
	.clk(clk),
	.d(\fp_functions_0|add_5~9_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][56]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][56] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][56] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][57] (
	.clk(clk),
	.d(\fp_functions_0|add_5~13_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][57]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][57] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][57] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][58] (
	.clk(clk),
	.d(\fp_functions_0|add_5~17_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][58]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][58] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][58] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][59] (
	.clk(clk),
	.d(\fp_functions_0|add_5~21_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][59]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][59] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][59] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][60] (
	.clk(clk),
	.d(\fp_functions_0|add_5~25_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][60]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][60] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][60] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][61] (
	.clk(clk),
	.d(\fp_functions_0|add_5~29_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][61]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][61] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][61] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][62] (
	.clk(clk),
	.d(\fp_functions_0|add_5~33_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][62]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][62] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][62] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][63] (
	.clk(clk),
	.d(\fp_functions_0|add_5~37_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][63]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][63] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][63] .power_up = "low";

dffeas \fp_functions_0|redist14|delay_signals[3][0] (
	.clk(clk),
	.d(\fp_functions_0|redist14|delay_signals[4][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist14|delay_signals[3][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist14|delay_signals[3][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist14|delay_signals[3][0] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][0] (
	.clk(clk),
	.d(\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][0] .power_up = "low";

dffeas \fp_functions_0|roundBit_uid65_fpMulTest_delay|delay_signals[0][0] (
	.clk(clk),
	.d(\fp_functions_0|reduce_nor_7~combout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|roundBit_uid65_fpMulTest_delay|delay_signals[0][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|roundBit_uid65_fpMulTest_delay|delay_signals[0][0] .is_wysiwyg = "true";
defparam \fp_functions_0|roundBit_uid65_fpMulTest_delay|delay_signals[0][0] .power_up = "low";

dffeas \fp_functions_0|redist18|delay_signals[3][0] (
	.clk(clk),
	.d(\fp_functions_0|redist18|delay_signals[4][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist18|delay_signals[3][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist18|delay_signals[3][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist18|delay_signals[3][0] .power_up = "low";

dffeas \fp_functions_0|redist17|delay_signals[3][0] (
	.clk(clk),
	.d(\fp_functions_0|redist17|delay_signals[4][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist17|delay_signals[3][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist17|delay_signals[3][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist17|delay_signals[3][0] .power_up = "low";

dffeas \fp_functions_0|redist20|delay_signals[3][0] (
	.clk(clk),
	.d(\fp_functions_0|redist20|delay_signals[4][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist20|delay_signals[3][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist20|delay_signals[3][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist20|delay_signals[3][0] .power_up = "low";

dffeas \fp_functions_0|redist21|delay_signals[3][0] (
	.clk(clk),
	.d(\fp_functions_0|redist21|delay_signals[4][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist21|delay_signals[3][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist21|delay_signals[3][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist21|delay_signals[3][0] .power_up = "low";

dffeas \fp_functions_0|redist16|delay_signals[3][0] (
	.clk(clk),
	.d(\fp_functions_0|redist16|delay_signals[4][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist16|delay_signals[3][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist16|delay_signals[3][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist16|delay_signals[3][0] .power_up = "low";

dffeas \fp_functions_0|redist19|delay_signals[3][0] (
	.clk(clk),
	.d(\fp_functions_0|redist19|delay_signals[4][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist19|delay_signals[3][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist19|delay_signals[3][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist19|delay_signals[3][0] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][66] (
	.clk(clk),
	.d(\fp_functions_0|add_5~41_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][66]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][66] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][66] .power_up = "low";

dffeas \fp_functions_0|redist9|delay_signals[0][13] (
	.clk(clk),
	.d(\fp_functions_0|add_6~261_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist9|delay_signals[0][13]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist9|delay_signals[0][13] .is_wysiwyg = "true";
defparam \fp_functions_0|redist9|delay_signals[0][13] .power_up = "low";

dffeas \fp_functions_0|redist15_outputreg|delay_signals[0][0] (
	.clk(clk),
	.d(\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist15_outputreg|delay_signals[0][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist15_outputreg|delay_signals[0][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist15_outputreg|delay_signals[0][0] .power_up = "low";

dffeas \fp_functions_0|redist13|delay_signals[1][0] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][105]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist13|delay_signals[1][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist13|delay_signals[1][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist13|delay_signals[1][0] .power_up = "low";

dffeas \fp_functions_0|redist14|delay_signals[4][0] (
	.clk(clk),
	.d(\fp_functions_0|redist14|delay_signals[5][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist14|delay_signals[4][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist14|delay_signals[4][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist14|delay_signals[4][0] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][52] (
	.clk(clk),
	.d(\fp_functions_0|add_1~1_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][52]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][52] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][52] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][53] (
	.clk(clk),
	.d(\fp_functions_0|add_1~5_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][53]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][53] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][53] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][105] (
	.clk(clk),
	.d(\fp_functions_0|add_1~9_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][105]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][105] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][105] .power_up = "low";

dffeas \fp_functions_0|redist12|delay_signals[0][48] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][48]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist12|delay_signals[0][48]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist12|delay_signals[0][48] .is_wysiwyg = "true";
defparam \fp_functions_0|redist12|delay_signals[0][48] .power_up = "low";

dffeas \fp_functions_0|redist12|delay_signals[0][49] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][49]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist12|delay_signals[0][49]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist12|delay_signals[0][49] .is_wysiwyg = "true";
defparam \fp_functions_0|redist12|delay_signals[0][49] .power_up = "low";

dffeas \fp_functions_0|redist12|delay_signals[0][50] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][50]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist12|delay_signals[0][50]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist12|delay_signals[0][50] .is_wysiwyg = "true";
defparam \fp_functions_0|redist12|delay_signals[0][50] .power_up = "low";

dffeas \fp_functions_0|redist12|delay_signals[0][51] (
	.clk(clk),
	.d(\fp_functions_0|i5343~0_combout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist12|delay_signals[0][51]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist12|delay_signals[0][51] .is_wysiwyg = "true";
defparam \fp_functions_0|redist12|delay_signals[0][51] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|reduce_nor_7~0 (
	.dataa(!\fp_functions_0|redist12|delay_signals[0][48]~q ),
	.datab(!\fp_functions_0|redist12|delay_signals[0][49]~q ),
	.datac(!\fp_functions_0|redist12|delay_signals[0][50]~q ),
	.datad(!\fp_functions_0|redist12|delay_signals[0][51]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|reduce_nor_7~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|reduce_nor_7~0 .extended_lut = "off";
defparam \fp_functions_0|reduce_nor_7~0 .lut_mask = 64'h8000800080008000;
defparam \fp_functions_0|reduce_nor_7~0 .shared_arith = "off";

dffeas \fp_functions_0|redist12|delay_signals[0][41] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][41]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist12|delay_signals[0][41]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist12|delay_signals[0][41] .is_wysiwyg = "true";
defparam \fp_functions_0|redist12|delay_signals[0][41] .power_up = "low";

dffeas \fp_functions_0|redist12|delay_signals[0][46] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][46]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist12|delay_signals[0][46]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist12|delay_signals[0][46] .is_wysiwyg = "true";
defparam \fp_functions_0|redist12|delay_signals[0][46] .power_up = "low";

dffeas \fp_functions_0|redist12|delay_signals[0][47] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][47]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist12|delay_signals[0][47]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist12|delay_signals[0][47] .is_wysiwyg = "true";
defparam \fp_functions_0|redist12|delay_signals[0][47] .power_up = "low";

dffeas \fp_functions_0|redist12|delay_signals[0][42] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][42]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist12|delay_signals[0][42]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist12|delay_signals[0][42] .is_wysiwyg = "true";
defparam \fp_functions_0|redist12|delay_signals[0][42] .power_up = "low";

dffeas \fp_functions_0|redist12|delay_signals[0][43] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][43]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist12|delay_signals[0][43]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist12|delay_signals[0][43] .is_wysiwyg = "true";
defparam \fp_functions_0|redist12|delay_signals[0][43] .power_up = "low";

dffeas \fp_functions_0|redist12|delay_signals[0][44] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][44]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist12|delay_signals[0][44]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist12|delay_signals[0][44] .is_wysiwyg = "true";
defparam \fp_functions_0|redist12|delay_signals[0][44] .power_up = "low";

dffeas \fp_functions_0|redist12|delay_signals[0][45] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][45]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist12|delay_signals[0][45]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist12|delay_signals[0][45] .is_wysiwyg = "true";
defparam \fp_functions_0|redist12|delay_signals[0][45] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|reduce_nor_7~1 (
	.dataa(!\fp_functions_0|redist12|delay_signals[0][42]~q ),
	.datab(!\fp_functions_0|redist12|delay_signals[0][43]~q ),
	.datac(!\fp_functions_0|redist12|delay_signals[0][44]~q ),
	.datad(!\fp_functions_0|redist12|delay_signals[0][45]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|reduce_nor_7~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|reduce_nor_7~1 .extended_lut = "off";
defparam \fp_functions_0|reduce_nor_7~1 .lut_mask = 64'h8000800080008000;
defparam \fp_functions_0|reduce_nor_7~1 .shared_arith = "off";

dffeas \fp_functions_0|redist12|delay_signals[0][36] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][36]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist12|delay_signals[0][36]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist12|delay_signals[0][36] .is_wysiwyg = "true";
defparam \fp_functions_0|redist12|delay_signals[0][36] .power_up = "low";

dffeas \fp_functions_0|redist12|delay_signals[0][37] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][37]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist12|delay_signals[0][37]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist12|delay_signals[0][37] .is_wysiwyg = "true";
defparam \fp_functions_0|redist12|delay_signals[0][37] .power_up = "low";

dffeas \fp_functions_0|redist12|delay_signals[0][38] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][38]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist12|delay_signals[0][38]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist12|delay_signals[0][38] .is_wysiwyg = "true";
defparam \fp_functions_0|redist12|delay_signals[0][38] .power_up = "low";

dffeas \fp_functions_0|redist12|delay_signals[0][39] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][39]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist12|delay_signals[0][39]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist12|delay_signals[0][39] .is_wysiwyg = "true";
defparam \fp_functions_0|redist12|delay_signals[0][39] .power_up = "low";

dffeas \fp_functions_0|redist12|delay_signals[0][40] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][40]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist12|delay_signals[0][40]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist12|delay_signals[0][40] .is_wysiwyg = "true";
defparam \fp_functions_0|redist12|delay_signals[0][40] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|reduce_nor_7~2 (
	.dataa(!\fp_functions_0|redist12|delay_signals[0][36]~q ),
	.datab(!\fp_functions_0|redist12|delay_signals[0][37]~q ),
	.datac(!\fp_functions_0|redist12|delay_signals[0][38]~q ),
	.datad(!\fp_functions_0|redist12|delay_signals[0][39]~q ),
	.datae(!\fp_functions_0|redist12|delay_signals[0][40]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|reduce_nor_7~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|reduce_nor_7~2 .extended_lut = "off";
defparam \fp_functions_0|reduce_nor_7~2 .lut_mask = 64'h8000000080000000;
defparam \fp_functions_0|reduce_nor_7~2 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|reduce_nor_7~3 (
	.dataa(!\fp_functions_0|redist12|delay_signals[0][41]~q ),
	.datab(!\fp_functions_0|redist12|delay_signals[0][46]~q ),
	.datac(!\fp_functions_0|redist12|delay_signals[0][47]~q ),
	.datad(!\fp_functions_0|reduce_nor_7~1_combout ),
	.datae(!\fp_functions_0|reduce_nor_7~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|reduce_nor_7~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|reduce_nor_7~3 .extended_lut = "off";
defparam \fp_functions_0|reduce_nor_7~3 .lut_mask = 64'h0000008000000080;
defparam \fp_functions_0|reduce_nor_7~3 .shared_arith = "off";

dffeas \fp_functions_0|redist12|delay_signals[0][29] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][29]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist12|delay_signals[0][29]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist12|delay_signals[0][29] .is_wysiwyg = "true";
defparam \fp_functions_0|redist12|delay_signals[0][29] .power_up = "low";

dffeas \fp_functions_0|redist12|delay_signals[0][35] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][35]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist12|delay_signals[0][35]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist12|delay_signals[0][35] .is_wysiwyg = "true";
defparam \fp_functions_0|redist12|delay_signals[0][35] .power_up = "low";

dffeas \fp_functions_0|redist12|delay_signals[0][24] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][24]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist12|delay_signals[0][24]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist12|delay_signals[0][24] .is_wysiwyg = "true";
defparam \fp_functions_0|redist12|delay_signals[0][24] .power_up = "low";

dffeas \fp_functions_0|redist12|delay_signals[0][25] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][25]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist12|delay_signals[0][25]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist12|delay_signals[0][25] .is_wysiwyg = "true";
defparam \fp_functions_0|redist12|delay_signals[0][25] .power_up = "low";

dffeas \fp_functions_0|redist12|delay_signals[0][26] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][26]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist12|delay_signals[0][26]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist12|delay_signals[0][26] .is_wysiwyg = "true";
defparam \fp_functions_0|redist12|delay_signals[0][26] .power_up = "low";

dffeas \fp_functions_0|redist12|delay_signals[0][27] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][27]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist12|delay_signals[0][27]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist12|delay_signals[0][27] .is_wysiwyg = "true";
defparam \fp_functions_0|redist12|delay_signals[0][27] .power_up = "low";

dffeas \fp_functions_0|redist12|delay_signals[0][28] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][28]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist12|delay_signals[0][28]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist12|delay_signals[0][28] .is_wysiwyg = "true";
defparam \fp_functions_0|redist12|delay_signals[0][28] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|reduce_nor_7~4 (
	.dataa(!\fp_functions_0|redist12|delay_signals[0][24]~q ),
	.datab(!\fp_functions_0|redist12|delay_signals[0][25]~q ),
	.datac(!\fp_functions_0|redist12|delay_signals[0][26]~q ),
	.datad(!\fp_functions_0|redist12|delay_signals[0][27]~q ),
	.datae(!\fp_functions_0|redist12|delay_signals[0][28]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|reduce_nor_7~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|reduce_nor_7~4 .extended_lut = "off";
defparam \fp_functions_0|reduce_nor_7~4 .lut_mask = 64'h8000000080000000;
defparam \fp_functions_0|reduce_nor_7~4 .shared_arith = "off";

dffeas \fp_functions_0|redist12|delay_signals[0][30] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][30]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist12|delay_signals[0][30]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist12|delay_signals[0][30] .is_wysiwyg = "true";
defparam \fp_functions_0|redist12|delay_signals[0][30] .power_up = "low";

dffeas \fp_functions_0|redist12|delay_signals[0][31] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][31]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist12|delay_signals[0][31]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist12|delay_signals[0][31] .is_wysiwyg = "true";
defparam \fp_functions_0|redist12|delay_signals[0][31] .power_up = "low";

dffeas \fp_functions_0|redist12|delay_signals[0][32] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][32]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist12|delay_signals[0][32]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist12|delay_signals[0][32] .is_wysiwyg = "true";
defparam \fp_functions_0|redist12|delay_signals[0][32] .power_up = "low";

dffeas \fp_functions_0|redist12|delay_signals[0][33] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][33]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist12|delay_signals[0][33]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist12|delay_signals[0][33] .is_wysiwyg = "true";
defparam \fp_functions_0|redist12|delay_signals[0][33] .power_up = "low";

dffeas \fp_functions_0|redist12|delay_signals[0][34] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][34]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist12|delay_signals[0][34]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist12|delay_signals[0][34] .is_wysiwyg = "true";
defparam \fp_functions_0|redist12|delay_signals[0][34] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|reduce_nor_7~5 (
	.dataa(!\fp_functions_0|redist12|delay_signals[0][30]~q ),
	.datab(!\fp_functions_0|redist12|delay_signals[0][31]~q ),
	.datac(!\fp_functions_0|redist12|delay_signals[0][32]~q ),
	.datad(!\fp_functions_0|redist12|delay_signals[0][33]~q ),
	.datae(!\fp_functions_0|redist12|delay_signals[0][34]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|reduce_nor_7~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|reduce_nor_7~5 .extended_lut = "off";
defparam \fp_functions_0|reduce_nor_7~5 .lut_mask = 64'h8000000080000000;
defparam \fp_functions_0|reduce_nor_7~5 .shared_arith = "off";

dffeas \fp_functions_0|redist12|delay_signals[0][17] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][17]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist12|delay_signals[0][17]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist12|delay_signals[0][17] .is_wysiwyg = "true";
defparam \fp_functions_0|redist12|delay_signals[0][17] .power_up = "low";

dffeas \fp_functions_0|redist12|delay_signals[0][23] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][23]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist12|delay_signals[0][23]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist12|delay_signals[0][23] .is_wysiwyg = "true";
defparam \fp_functions_0|redist12|delay_signals[0][23] .power_up = "low";

dffeas \fp_functions_0|redist12|delay_signals[0][12] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][12]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist12|delay_signals[0][12]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist12|delay_signals[0][12] .is_wysiwyg = "true";
defparam \fp_functions_0|redist12|delay_signals[0][12] .power_up = "low";

dffeas \fp_functions_0|redist12|delay_signals[0][13] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][13]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist12|delay_signals[0][13]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist12|delay_signals[0][13] .is_wysiwyg = "true";
defparam \fp_functions_0|redist12|delay_signals[0][13] .power_up = "low";

dffeas \fp_functions_0|redist12|delay_signals[0][14] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][14]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist12|delay_signals[0][14]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist12|delay_signals[0][14] .is_wysiwyg = "true";
defparam \fp_functions_0|redist12|delay_signals[0][14] .power_up = "low";

dffeas \fp_functions_0|redist12|delay_signals[0][15] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][15]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist12|delay_signals[0][15]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist12|delay_signals[0][15] .is_wysiwyg = "true";
defparam \fp_functions_0|redist12|delay_signals[0][15] .power_up = "low";

dffeas \fp_functions_0|redist12|delay_signals[0][16] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][16]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist12|delay_signals[0][16]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist12|delay_signals[0][16] .is_wysiwyg = "true";
defparam \fp_functions_0|redist12|delay_signals[0][16] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|reduce_nor_7~6 (
	.dataa(!\fp_functions_0|redist12|delay_signals[0][12]~q ),
	.datab(!\fp_functions_0|redist12|delay_signals[0][13]~q ),
	.datac(!\fp_functions_0|redist12|delay_signals[0][14]~q ),
	.datad(!\fp_functions_0|redist12|delay_signals[0][15]~q ),
	.datae(!\fp_functions_0|redist12|delay_signals[0][16]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|reduce_nor_7~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|reduce_nor_7~6 .extended_lut = "off";
defparam \fp_functions_0|reduce_nor_7~6 .lut_mask = 64'h8000000080000000;
defparam \fp_functions_0|reduce_nor_7~6 .shared_arith = "off";

dffeas \fp_functions_0|redist12|delay_signals[0][18] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][18]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist12|delay_signals[0][18]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist12|delay_signals[0][18] .is_wysiwyg = "true";
defparam \fp_functions_0|redist12|delay_signals[0][18] .power_up = "low";

dffeas \fp_functions_0|redist12|delay_signals[0][19] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][19]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist12|delay_signals[0][19]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist12|delay_signals[0][19] .is_wysiwyg = "true";
defparam \fp_functions_0|redist12|delay_signals[0][19] .power_up = "low";

dffeas \fp_functions_0|redist12|delay_signals[0][20] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][20]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist12|delay_signals[0][20]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist12|delay_signals[0][20] .is_wysiwyg = "true";
defparam \fp_functions_0|redist12|delay_signals[0][20] .power_up = "low";

dffeas \fp_functions_0|redist12|delay_signals[0][21] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][21]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist12|delay_signals[0][21]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist12|delay_signals[0][21] .is_wysiwyg = "true";
defparam \fp_functions_0|redist12|delay_signals[0][21] .power_up = "low";

dffeas \fp_functions_0|redist12|delay_signals[0][22] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][22]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist12|delay_signals[0][22]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist12|delay_signals[0][22] .is_wysiwyg = "true";
defparam \fp_functions_0|redist12|delay_signals[0][22] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|reduce_nor_7~7 (
	.dataa(!\fp_functions_0|redist12|delay_signals[0][18]~q ),
	.datab(!\fp_functions_0|redist12|delay_signals[0][19]~q ),
	.datac(!\fp_functions_0|redist12|delay_signals[0][20]~q ),
	.datad(!\fp_functions_0|redist12|delay_signals[0][21]~q ),
	.datae(!\fp_functions_0|redist12|delay_signals[0][22]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|reduce_nor_7~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|reduce_nor_7~7 .extended_lut = "off";
defparam \fp_functions_0|reduce_nor_7~7 .lut_mask = 64'h8000000080000000;
defparam \fp_functions_0|reduce_nor_7~7 .shared_arith = "off";

dffeas \fp_functions_0|redist12|delay_signals[0][5] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][5]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist12|delay_signals[0][5]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist12|delay_signals[0][5] .is_wysiwyg = "true";
defparam \fp_functions_0|redist12|delay_signals[0][5] .power_up = "low";

dffeas \fp_functions_0|redist12|delay_signals[0][10] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][10]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist12|delay_signals[0][10]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist12|delay_signals[0][10] .is_wysiwyg = "true";
defparam \fp_functions_0|redist12|delay_signals[0][10] .power_up = "low";

dffeas \fp_functions_0|redist12|delay_signals[0][11] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][11]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist12|delay_signals[0][11]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist12|delay_signals[0][11] .is_wysiwyg = "true";
defparam \fp_functions_0|redist12|delay_signals[0][11] .power_up = "low";

dffeas \fp_functions_0|redist12|delay_signals[0][6] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][6]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist12|delay_signals[0][6]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist12|delay_signals[0][6] .is_wysiwyg = "true";
defparam \fp_functions_0|redist12|delay_signals[0][6] .power_up = "low";

dffeas \fp_functions_0|redist12|delay_signals[0][7] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][7]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist12|delay_signals[0][7]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist12|delay_signals[0][7] .is_wysiwyg = "true";
defparam \fp_functions_0|redist12|delay_signals[0][7] .power_up = "low";

dffeas \fp_functions_0|redist12|delay_signals[0][8] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][8]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist12|delay_signals[0][8]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist12|delay_signals[0][8] .is_wysiwyg = "true";
defparam \fp_functions_0|redist12|delay_signals[0][8] .power_up = "low";

dffeas \fp_functions_0|redist12|delay_signals[0][9] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][9]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist12|delay_signals[0][9]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist12|delay_signals[0][9] .is_wysiwyg = "true";
defparam \fp_functions_0|redist12|delay_signals[0][9] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|reduce_nor_7~8 (
	.dataa(!\fp_functions_0|redist12|delay_signals[0][6]~q ),
	.datab(!\fp_functions_0|redist12|delay_signals[0][7]~q ),
	.datac(!\fp_functions_0|redist12|delay_signals[0][8]~q ),
	.datad(!\fp_functions_0|redist12|delay_signals[0][9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|reduce_nor_7~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|reduce_nor_7~8 .extended_lut = "off";
defparam \fp_functions_0|reduce_nor_7~8 .lut_mask = 64'h8000800080008000;
defparam \fp_functions_0|reduce_nor_7~8 .shared_arith = "off";

dffeas \fp_functions_0|redist12|delay_signals[0][0] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist12|delay_signals[0][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist12|delay_signals[0][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist12|delay_signals[0][0] .power_up = "low";

dffeas \fp_functions_0|redist12|delay_signals[0][1] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][1]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist12|delay_signals[0][1]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist12|delay_signals[0][1] .is_wysiwyg = "true";
defparam \fp_functions_0|redist12|delay_signals[0][1] .power_up = "low";

dffeas \fp_functions_0|redist12|delay_signals[0][2] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][2]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist12|delay_signals[0][2]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist12|delay_signals[0][2] .is_wysiwyg = "true";
defparam \fp_functions_0|redist12|delay_signals[0][2] .power_up = "low";

dffeas \fp_functions_0|redist12|delay_signals[0][3] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][3]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist12|delay_signals[0][3]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist12|delay_signals[0][3] .is_wysiwyg = "true";
defparam \fp_functions_0|redist12|delay_signals[0][3] .power_up = "low";

dffeas \fp_functions_0|redist12|delay_signals[0][4] (
	.clk(clk),
	.d(\fp_functions_0|redist1|delay_signals[0][4]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist12|delay_signals[0][4]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist12|delay_signals[0][4] .is_wysiwyg = "true";
defparam \fp_functions_0|redist12|delay_signals[0][4] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|reduce_nor_7~9 (
	.dataa(!\fp_functions_0|redist12|delay_signals[0][0]~q ),
	.datab(!\fp_functions_0|redist12|delay_signals[0][1]~q ),
	.datac(!\fp_functions_0|redist12|delay_signals[0][2]~q ),
	.datad(!\fp_functions_0|redist12|delay_signals[0][3]~q ),
	.datae(!\fp_functions_0|redist12|delay_signals[0][4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|reduce_nor_7~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|reduce_nor_7~9 .extended_lut = "off";
defparam \fp_functions_0|reduce_nor_7~9 .lut_mask = 64'h8000000080000000;
defparam \fp_functions_0|reduce_nor_7~9 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|reduce_nor_7~10 (
	.dataa(!\fp_functions_0|redist12|delay_signals[0][5]~q ),
	.datab(!\fp_functions_0|redist12|delay_signals[0][10]~q ),
	.datac(!\fp_functions_0|redist12|delay_signals[0][11]~q ),
	.datad(!\fp_functions_0|reduce_nor_7~8_combout ),
	.datae(!\fp_functions_0|reduce_nor_7~9_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|reduce_nor_7~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|reduce_nor_7~10 .extended_lut = "off";
defparam \fp_functions_0|reduce_nor_7~10 .lut_mask = 64'h0000008000000080;
defparam \fp_functions_0|reduce_nor_7~10 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|reduce_nor_7 (
	.dataa(!\fp_functions_0|reduce_nor_7~0_combout ),
	.datab(!\fp_functions_0|reduce_nor_7~3_combout ),
	.datac(!\fp_functions_0|reduce_nor_7~4_combout ),
	.datad(!\fp_functions_0|reduce_nor_7~10_combout ),
	.datae(!\fp_functions_0|reduce_nor_7~11_combout ),
	.dataf(!\fp_functions_0|reduce_nor_7~12_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|reduce_nor_7~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|reduce_nor_7 .extended_lut = "off";
defparam \fp_functions_0|reduce_nor_7 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \fp_functions_0|reduce_nor_7 .shared_arith = "off";

dffeas \fp_functions_0|redist18|delay_signals[4][0] (
	.clk(clk),
	.d(\fp_functions_0|redist18|delay_signals[5][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist18|delay_signals[4][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist18|delay_signals[4][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist18|delay_signals[4][0] .power_up = "low";

dffeas \fp_functions_0|redist17|delay_signals[4][0] (
	.clk(clk),
	.d(\fp_functions_0|redist17|delay_signals[5][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist17|delay_signals[4][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist17|delay_signals[4][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist17|delay_signals[4][0] .power_up = "low";

dffeas \fp_functions_0|redist20|delay_signals[4][0] (
	.clk(clk),
	.d(\fp_functions_0|redist20|delay_signals[5][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist20|delay_signals[4][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist20|delay_signals[4][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist20|delay_signals[4][0] .power_up = "low";

dffeas \fp_functions_0|redist21|delay_signals[4][0] (
	.clk(clk),
	.d(\fp_functions_0|redist21|delay_signals[5][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist21|delay_signals[4][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist21|delay_signals[4][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist21|delay_signals[4][0] .power_up = "low";

dffeas \fp_functions_0|redist16|delay_signals[4][0] (
	.clk(clk),
	.d(\fp_functions_0|redist16|delay_signals[5][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist16|delay_signals[4][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist16|delay_signals[4][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist16|delay_signals[4][0] .power_up = "low";

dffeas \fp_functions_0|redist19|delay_signals[4][0] (
	.clk(clk),
	.d(\fp_functions_0|redist19|delay_signals[5][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist19|delay_signals[4][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist19|delay_signals[4][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist19|delay_signals[4][0] .power_up = "low";

dffeas \fp_functions_0|redist9|delay_signals[0][12] (
	.clk(clk),
	.d(\fp_functions_0|add_6~265_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist9|delay_signals[0][12]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist9|delay_signals[0][12] .is_wysiwyg = "true";
defparam \fp_functions_0|redist9|delay_signals[0][12] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][54] (
	.clk(clk),
	.d(\fp_functions_0|add_1~13_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][54]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][54] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][54] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][55] (
	.clk(clk),
	.d(\fp_functions_0|add_1~17_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][55]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][55] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][55] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][56] (
	.clk(clk),
	.d(\fp_functions_0|add_1~21_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][56]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][56] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][56] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][57] (
	.clk(clk),
	.d(\fp_functions_0|add_1~25_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][57]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][57] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][57] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][58] (
	.clk(clk),
	.d(\fp_functions_0|add_1~29_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][58]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][58] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][58] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][59] (
	.clk(clk),
	.d(\fp_functions_0|add_1~33_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][59]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][59] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][59] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][60] (
	.clk(clk),
	.d(\fp_functions_0|add_1~37_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][60]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][60] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][60] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][61] (
	.clk(clk),
	.d(\fp_functions_0|add_1~41_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][61]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][61] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][61] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][62] (
	.clk(clk),
	.d(\fp_functions_0|add_1~45_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][62]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][62] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][62] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][63] (
	.clk(clk),
	.d(\fp_functions_0|add_1~49_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][63]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][63] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][63] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][64] (
	.clk(clk),
	.d(\fp_functions_0|add_1~53_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][64]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][64] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][64] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][65] (
	.clk(clk),
	.d(\fp_functions_0|add_1~57_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][65]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][65] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][65] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][66] (
	.clk(clk),
	.d(\fp_functions_0|add_1~61_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][66]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][66] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][66] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][67] (
	.clk(clk),
	.d(\fp_functions_0|add_1~65_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][67]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][67] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][67] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][68] (
	.clk(clk),
	.d(\fp_functions_0|add_1~69_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][68]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][68] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][68] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][69] (
	.clk(clk),
	.d(\fp_functions_0|add_1~73_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][69]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][69] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][69] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][70] (
	.clk(clk),
	.d(\fp_functions_0|add_1~77_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][70]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][70] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][70] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][71] (
	.clk(clk),
	.d(\fp_functions_0|add_1~81_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][71]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][71] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][71] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][72] (
	.clk(clk),
	.d(\fp_functions_0|add_1~85_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][72]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][72] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][72] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][73] (
	.clk(clk),
	.d(\fp_functions_0|add_1~89_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][73]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][73] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][73] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][74] (
	.clk(clk),
	.d(\fp_functions_0|add_1~93_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][74]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][74] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][74] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][75] (
	.clk(clk),
	.d(\fp_functions_0|add_1~97_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][75]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][75] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][75] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][76] (
	.clk(clk),
	.d(\fp_functions_0|add_1~101_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][76]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][76] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][76] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][77] (
	.clk(clk),
	.d(\fp_functions_0|add_1~105_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][77]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][77] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][77] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][78] (
	.clk(clk),
	.d(\fp_functions_0|add_1~109_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][78]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][78] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][78] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][79] (
	.clk(clk),
	.d(\fp_functions_0|add_1~113_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][79]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][79] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][79] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][80] (
	.clk(clk),
	.d(\fp_functions_0|add_1~117_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][80]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][80] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][80] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][81] (
	.clk(clk),
	.d(\fp_functions_0|add_1~121_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][81]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][81] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][81] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][82] (
	.clk(clk),
	.d(\fp_functions_0|add_1~125_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][82]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][82] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][82] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][83] (
	.clk(clk),
	.d(\fp_functions_0|add_1~129_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][83]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][83] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][83] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][84] (
	.clk(clk),
	.d(\fp_functions_0|add_1~133_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][84]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][84] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][84] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][85] (
	.clk(clk),
	.d(\fp_functions_0|add_1~137_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][85]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][85] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][85] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][86] (
	.clk(clk),
	.d(\fp_functions_0|add_1~141_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][86]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][86] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][86] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][87] (
	.clk(clk),
	.d(\fp_functions_0|add_1~145_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][87]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][87] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][87] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][88] (
	.clk(clk),
	.d(\fp_functions_0|add_1~149_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][88]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][88] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][88] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][89] (
	.clk(clk),
	.d(\fp_functions_0|add_1~153_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][89]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][89] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][89] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][90] (
	.clk(clk),
	.d(\fp_functions_0|add_1~157_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][90]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][90] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][90] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][91] (
	.clk(clk),
	.d(\fp_functions_0|add_1~161_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][91]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][91] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][91] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][92] (
	.clk(clk),
	.d(\fp_functions_0|add_1~165_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][92]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][92] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][92] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][93] (
	.clk(clk),
	.d(\fp_functions_0|add_1~169_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][93]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][93] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][93] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][94] (
	.clk(clk),
	.d(\fp_functions_0|add_1~173_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][94]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][94] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][94] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][95] (
	.clk(clk),
	.d(\fp_functions_0|add_1~177_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][95]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][95] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][95] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][96] (
	.clk(clk),
	.d(\fp_functions_0|add_1~181_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][96]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][96] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][96] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][97] (
	.clk(clk),
	.d(\fp_functions_0|add_1~185_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][97]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][97] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][97] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][98] (
	.clk(clk),
	.d(\fp_functions_0|add_1~189_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][98]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][98] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][98] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][99] (
	.clk(clk),
	.d(\fp_functions_0|add_1~193_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][99]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][99] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][99] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][100] (
	.clk(clk),
	.d(\fp_functions_0|add_1~197_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][100]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][100] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][100] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][101] (
	.clk(clk),
	.d(\fp_functions_0|add_1~201_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][101]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][101] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][101] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][102] (
	.clk(clk),
	.d(\fp_functions_0|add_1~205_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][102]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][102] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][102] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][103] (
	.clk(clk),
	.d(\fp_functions_0|add_1~209_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][103]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][103] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][103] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][104] (
	.clk(clk),
	.d(\fp_functions_0|add_1~213_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][104]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][104] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][104] .power_up = "low";

dffeas \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[0] (
	.clk(clk),
	.d(\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_wire[0] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\fp_functions_0|i5762~combout ),
	.q(\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[0] .power_up = "low";

dffeas \fp_functions_0|redist15_outputreg|delay_signals[0][1] (
	.clk(clk),
	.d(\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[1]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist15_outputreg|delay_signals[0][1]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist15_outputreg|delay_signals[0][1] .is_wysiwyg = "true";
defparam \fp_functions_0|redist15_outputreg|delay_signals[0][1] .power_up = "low";

dffeas \fp_functions_0|redist15_outputreg|delay_signals[0][2] (
	.clk(clk),
	.d(\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[2]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist15_outputreg|delay_signals[0][2]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist15_outputreg|delay_signals[0][2] .is_wysiwyg = "true";
defparam \fp_functions_0|redist15_outputreg|delay_signals[0][2] .power_up = "low";

dffeas \fp_functions_0|redist15_outputreg|delay_signals[0][3] (
	.clk(clk),
	.d(\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[3]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist15_outputreg|delay_signals[0][3]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist15_outputreg|delay_signals[0][3] .is_wysiwyg = "true";
defparam \fp_functions_0|redist15_outputreg|delay_signals[0][3] .power_up = "low";

dffeas \fp_functions_0|redist15_outputreg|delay_signals[0][4] (
	.clk(clk),
	.d(\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[4]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist15_outputreg|delay_signals[0][4]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist15_outputreg|delay_signals[0][4] .is_wysiwyg = "true";
defparam \fp_functions_0|redist15_outputreg|delay_signals[0][4] .power_up = "low";

dffeas \fp_functions_0|redist15_outputreg|delay_signals[0][5] (
	.clk(clk),
	.d(\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[5]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist15_outputreg|delay_signals[0][5]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist15_outputreg|delay_signals[0][5] .is_wysiwyg = "true";
defparam \fp_functions_0|redist15_outputreg|delay_signals[0][5] .power_up = "low";

dffeas \fp_functions_0|redist15_outputreg|delay_signals[0][6] (
	.clk(clk),
	.d(\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[6]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist15_outputreg|delay_signals[0][6]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist15_outputreg|delay_signals[0][6] .is_wysiwyg = "true";
defparam \fp_functions_0|redist15_outputreg|delay_signals[0][6] .power_up = "low";

dffeas \fp_functions_0|redist15_outputreg|delay_signals[0][7] (
	.clk(clk),
	.d(\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[7]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist15_outputreg|delay_signals[0][7]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist15_outputreg|delay_signals[0][7] .is_wysiwyg = "true";
defparam \fp_functions_0|redist15_outputreg|delay_signals[0][7] .power_up = "low";

dffeas \fp_functions_0|redist15_outputreg|delay_signals[0][8] (
	.clk(clk),
	.d(\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[8]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist15_outputreg|delay_signals[0][8]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist15_outputreg|delay_signals[0][8] .is_wysiwyg = "true";
defparam \fp_functions_0|redist15_outputreg|delay_signals[0][8] .power_up = "low";

dffeas \fp_functions_0|redist15_outputreg|delay_signals[0][9] (
	.clk(clk),
	.d(\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[9]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist15_outputreg|delay_signals[0][9]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist15_outputreg|delay_signals[0][9] .is_wysiwyg = "true";
defparam \fp_functions_0|redist15_outputreg|delay_signals[0][9] .power_up = "low";

dffeas \fp_functions_0|redist15_outputreg|delay_signals[0][10] (
	.clk(clk),
	.d(\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[10]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist15_outputreg|delay_signals[0][10]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist15_outputreg|delay_signals[0][10] .is_wysiwyg = "true";
defparam \fp_functions_0|redist15_outputreg|delay_signals[0][10] .power_up = "low";

dffeas \fp_functions_0|redist14|delay_signals[5][0] (
	.clk(clk),
	.d(\fp_functions_0|redist14|delay_signals[6][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist14|delay_signals[5][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist14|delay_signals[5][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist14|delay_signals[5][0] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][51] (
	.clk(clk),
	.d(\fp_functions_0|add_1~217_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][51]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][51] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][51] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][48] (
	.clk(clk),
	.d(\fp_functions_0|add_1~221_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][48]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][48] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][48] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][49] (
	.clk(clk),
	.d(\fp_functions_0|add_1~225_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][49]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][49] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][49] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][50] (
	.clk(clk),
	.d(\fp_functions_0|add_1~229_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][50]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][50] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][50] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|i5343~0 (
	.dataa(!\fp_functions_0|redist1|delay_signals[0][105]~q ),
	.datab(!\fp_functions_0|redist1|delay_signals[0][51]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|i5343~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|i5343~0 .extended_lut = "off";
defparam \fp_functions_0|i5343~0 .lut_mask = 64'h1111111111111111;
defparam \fp_functions_0|i5343~0 .shared_arith = "off";

dffeas \fp_functions_0|redist1|delay_signals[0][41] (
	.clk(clk),
	.d(\fp_functions_0|add_1~233_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][41]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][41] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][41] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][46] (
	.clk(clk),
	.d(\fp_functions_0|add_1~237_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][46]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][46] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][46] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][47] (
	.clk(clk),
	.d(\fp_functions_0|add_1~241_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][47]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][47] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][47] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][42] (
	.clk(clk),
	.d(\fp_functions_0|add_1~245_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][42]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][42] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][42] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][43] (
	.clk(clk),
	.d(\fp_functions_0|add_1~249_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][43]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][43] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][43] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][44] (
	.clk(clk),
	.d(\fp_functions_0|add_1~253_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][44]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][44] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][44] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][45] (
	.clk(clk),
	.d(\fp_functions_0|add_1~257_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][45]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][45] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][45] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][36] (
	.clk(clk),
	.d(\fp_functions_0|add_1~261_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][36]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][36] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][36] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][37] (
	.clk(clk),
	.d(\fp_functions_0|add_1~265_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][37]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][37] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][37] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][38] (
	.clk(clk),
	.d(\fp_functions_0|add_1~269_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][38]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][38] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][38] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][39] (
	.clk(clk),
	.d(\fp_functions_0|add_1~273_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][39]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][39] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][39] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][40] (
	.clk(clk),
	.d(\fp_functions_0|add_1~277_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][40]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][40] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][40] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][29] (
	.clk(clk),
	.d(\fp_functions_0|add_1~281_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][29]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][29] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][29] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][35] (
	.clk(clk),
	.d(\fp_functions_0|add_1~285_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][35]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][35] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][35] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][24] (
	.clk(clk),
	.d(\fp_functions_0|redist3|delay_signals[0][26]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][24]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][24] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][24] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][25] (
	.clk(clk),
	.d(\fp_functions_0|add_1~289_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][25]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][25] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][25] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][26] (
	.clk(clk),
	.d(\fp_functions_0|add_1~293_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][26]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][26] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][26] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][27] (
	.clk(clk),
	.d(\fp_functions_0|add_1~297_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][27]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][27] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][27] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][28] (
	.clk(clk),
	.d(\fp_functions_0|add_1~301_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][28]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][28] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][28] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][30] (
	.clk(clk),
	.d(\fp_functions_0|add_1~305_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][30]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][30] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][30] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][31] (
	.clk(clk),
	.d(\fp_functions_0|add_1~309_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][31]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][31] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][31] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][32] (
	.clk(clk),
	.d(\fp_functions_0|add_1~313_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][32]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][32] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][32] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][33] (
	.clk(clk),
	.d(\fp_functions_0|add_1~317_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][33]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][33] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][33] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][34] (
	.clk(clk),
	.d(\fp_functions_0|add_1~321_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][34]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][34] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][34] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][17] (
	.clk(clk),
	.d(\fp_functions_0|redist3|delay_signals[0][19]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][17]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][17] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][17] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][23] (
	.clk(clk),
	.d(\fp_functions_0|redist3|delay_signals[0][25]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][23]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][23] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][23] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][12] (
	.clk(clk),
	.d(\fp_functions_0|redist3|delay_signals[0][14]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][12]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][12] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][12] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][13] (
	.clk(clk),
	.d(\fp_functions_0|redist3|delay_signals[0][15]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][13]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][13] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][13] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][14] (
	.clk(clk),
	.d(\fp_functions_0|redist3|delay_signals[0][16]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][14]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][14] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][14] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][15] (
	.clk(clk),
	.d(\fp_functions_0|redist3|delay_signals[0][17]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][15]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][15] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][15] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][16] (
	.clk(clk),
	.d(\fp_functions_0|redist3|delay_signals[0][18]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][16]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][16] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][16] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][18] (
	.clk(clk),
	.d(\fp_functions_0|redist3|delay_signals[0][20]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][18]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][18] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][18] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][19] (
	.clk(clk),
	.d(\fp_functions_0|redist3|delay_signals[0][21]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][19]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][19] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][19] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][20] (
	.clk(clk),
	.d(\fp_functions_0|redist3|delay_signals[0][22]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][20]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][20] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][20] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][21] (
	.clk(clk),
	.d(\fp_functions_0|redist3|delay_signals[0][23]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][21]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][21] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][21] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][22] (
	.clk(clk),
	.d(\fp_functions_0|redist3|delay_signals[0][24]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][22]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][22] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][22] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][5] (
	.clk(clk),
	.d(\fp_functions_0|redist3|delay_signals[0][7]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][5]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][5] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][5] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][10] (
	.clk(clk),
	.d(\fp_functions_0|redist3|delay_signals[0][12]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][10]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][10] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][10] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][11] (
	.clk(clk),
	.d(\fp_functions_0|redist3|delay_signals[0][13]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][11]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][11] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][11] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][6] (
	.clk(clk),
	.d(\fp_functions_0|redist3|delay_signals[0][8]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][6]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][6] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][6] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][7] (
	.clk(clk),
	.d(\fp_functions_0|redist3|delay_signals[0][9]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][7]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][7] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][7] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][8] (
	.clk(clk),
	.d(\fp_functions_0|redist3|delay_signals[0][10]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][8]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][8] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][8] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][9] (
	.clk(clk),
	.d(\fp_functions_0|redist3|delay_signals[0][11]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][9]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][9] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][9] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][0] (
	.clk(clk),
	.d(\fp_functions_0|redist3|delay_signals[0][2]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][0] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][1] (
	.clk(clk),
	.d(\fp_functions_0|redist3|delay_signals[0][3]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][1]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][1] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][1] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][2] (
	.clk(clk),
	.d(\fp_functions_0|redist3|delay_signals[0][4]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][2]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][2] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][2] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][3] (
	.clk(clk),
	.d(\fp_functions_0|redist3|delay_signals[0][5]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][3]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][3] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][3] .power_up = "low";

dffeas \fp_functions_0|redist1|delay_signals[0][4] (
	.clk(clk),
	.d(\fp_functions_0|redist3|delay_signals[0][6]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist1|delay_signals[0][4]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist1|delay_signals[0][4] .is_wysiwyg = "true";
defparam \fp_functions_0|redist1|delay_signals[0][4] .power_up = "low";

dffeas \fp_functions_0|redist18|delay_signals[5][0] (
	.clk(clk),
	.d(\fp_functions_0|redist18|delay_signals[6][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist18|delay_signals[5][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist18|delay_signals[5][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist18|delay_signals[5][0] .power_up = "low";

dffeas \fp_functions_0|redist17|delay_signals[5][0] (
	.clk(clk),
	.d(\fp_functions_0|redist17|delay_signals[6][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist17|delay_signals[5][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist17|delay_signals[5][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist17|delay_signals[5][0] .power_up = "low";

dffeas \fp_functions_0|redist20|delay_signals[5][0] (
	.clk(clk),
	.d(\fp_functions_0|redist20|delay_signals[6][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist20|delay_signals[5][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist20|delay_signals[5][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist20|delay_signals[5][0] .power_up = "low";

dffeas \fp_functions_0|redist21|delay_signals[5][0] (
	.clk(clk),
	.d(\fp_functions_0|redist21|delay_signals[6][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist21|delay_signals[5][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist21|delay_signals[5][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist21|delay_signals[5][0] .power_up = "low";

dffeas \fp_functions_0|redist16|delay_signals[5][0] (
	.clk(clk),
	.d(\fp_functions_0|redist16|delay_signals[6][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist16|delay_signals[5][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist16|delay_signals[5][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist16|delay_signals[5][0] .power_up = "low";

dffeas \fp_functions_0|redist19|delay_signals[5][0] (
	.clk(clk),
	.d(\fp_functions_0|redist19|delay_signals[6][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist19|delay_signals[5][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist19|delay_signals[5][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist19|delay_signals[5][0] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][65] (
	.clk(clk),
	.d(\fp_functions_0|add_5~45_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][65]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][65] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][65] .power_up = "low";

dffeas \fp_functions_0|redist9|delay_signals[0][11] (
	.clk(clk),
	.d(\fp_functions_0|add_6~269_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist9|delay_signals[0][11]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist9|delay_signals[0][11] .is_wysiwyg = "true";
defparam \fp_functions_0|redist9|delay_signals[0][11] .power_up = "low";

dffeas \fp_functions_0|redist15_sticky_ena_q[0] (
	.clk(clk),
	.d(\fp_functions_0|redist15_sticky_ena_q[0]~0_combout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\fp_functions_0|redist15_sticky_ena_q[0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist15_sticky_ena_q[0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist15_sticky_ena_q[0] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|i5762 (
	.dataa(!en[0]),
	.datab(!\fp_functions_0|redist15_sticky_ena_q[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|i5762~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|i5762 .extended_lut = "off";
defparam \fp_functions_0|i5762 .lut_mask = 64'h1111111111111111;
defparam \fp_functions_0|i5762 .shared_arith = "off";

dffeas \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[1] (
	.clk(clk),
	.d(\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_wire[1] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\fp_functions_0|i5762~combout ),
	.q(\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[1]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[1] .is_wysiwyg = "true";
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[1] .power_up = "low";

dffeas \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[2] (
	.clk(clk),
	.d(\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_wire[2] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\fp_functions_0|i5762~combout ),
	.q(\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[2]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[2] .is_wysiwyg = "true";
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[2] .power_up = "low";

dffeas \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[3] (
	.clk(clk),
	.d(\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_wire[3] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\fp_functions_0|i5762~combout ),
	.q(\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[3]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[3] .is_wysiwyg = "true";
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[3] .power_up = "low";

dffeas \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[4] (
	.clk(clk),
	.d(\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_wire[4] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\fp_functions_0|i5762~combout ),
	.q(\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[4]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[4] .is_wysiwyg = "true";
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[4] .power_up = "low";

dffeas \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[5] (
	.clk(clk),
	.d(\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_wire[5] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\fp_functions_0|i5762~combout ),
	.q(\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[5]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[5] .is_wysiwyg = "true";
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[5] .power_up = "low";

dffeas \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[6] (
	.clk(clk),
	.d(\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_wire[6] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\fp_functions_0|i5762~combout ),
	.q(\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[6]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[6] .is_wysiwyg = "true";
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[6] .power_up = "low";

dffeas \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[7] (
	.clk(clk),
	.d(\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_wire[7] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\fp_functions_0|i5762~combout ),
	.q(\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[7]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[7] .is_wysiwyg = "true";
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[7] .power_up = "low";

dffeas \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[8] (
	.clk(clk),
	.d(\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_wire[8] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\fp_functions_0|i5762~combout ),
	.q(\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[8]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[8] .is_wysiwyg = "true";
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[8] .power_up = "low";

dffeas \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[9] (
	.clk(clk),
	.d(\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_wire[9] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\fp_functions_0|i5762~combout ),
	.q(\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[9]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[9] .is_wysiwyg = "true";
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[9] .power_up = "low";

dffeas \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[10] (
	.clk(clk),
	.d(\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_wire[10] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\fp_functions_0|i5762~combout ),
	.q(\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[10]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[10] .is_wysiwyg = "true";
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[10] .power_up = "low";

dffeas \fp_functions_0|redist14|delay_signals[6][0] (
	.clk(clk),
	.d(\fp_functions_0|redist14|delay_signals[7][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist14|delay_signals[6][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist14|delay_signals[6][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist14|delay_signals[6][0] .power_up = "low";

dffeas \fp_functions_0|redist0|delay_signals[0][27] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][27]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist0|delay_signals[0][27]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist0|delay_signals[0][27] .is_wysiwyg = "true";
defparam \fp_functions_0|redist0|delay_signals[0][27] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][27] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][27]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][27] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][27] .power_up = "low";

dffeas \fp_functions_0|redist0|delay_signals[0][28] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][28]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist0|delay_signals[0][28]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist0|delay_signals[0][28] .is_wysiwyg = "true";
defparam \fp_functions_0|redist0|delay_signals[0][28] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][28] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][1]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][28]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][28] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][28] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][80] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][53]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][80]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][80] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][80] .power_up = "low";

dffeas \fp_functions_0|redist3|delay_signals[0][26] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][26]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist3|delay_signals[0][26]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist3|delay_signals[0][26] .is_wysiwyg = "true";
defparam \fp_functions_0|redist3|delay_signals[0][26] .power_up = "low";

dffeas \fp_functions_0|redist3|delay_signals[0][19] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][19]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist3|delay_signals[0][19]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist3|delay_signals[0][19] .is_wysiwyg = "true";
defparam \fp_functions_0|redist3|delay_signals[0][19] .power_up = "low";

dffeas \fp_functions_0|redist3|delay_signals[0][25] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][25]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist3|delay_signals[0][25]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist3|delay_signals[0][25] .is_wysiwyg = "true";
defparam \fp_functions_0|redist3|delay_signals[0][25] .power_up = "low";

dffeas \fp_functions_0|redist3|delay_signals[0][14] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][14]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist3|delay_signals[0][14]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist3|delay_signals[0][14] .is_wysiwyg = "true";
defparam \fp_functions_0|redist3|delay_signals[0][14] .power_up = "low";

dffeas \fp_functions_0|redist3|delay_signals[0][15] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][15]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist3|delay_signals[0][15]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist3|delay_signals[0][15] .is_wysiwyg = "true";
defparam \fp_functions_0|redist3|delay_signals[0][15] .power_up = "low";

dffeas \fp_functions_0|redist3|delay_signals[0][16] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][16]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist3|delay_signals[0][16]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist3|delay_signals[0][16] .is_wysiwyg = "true";
defparam \fp_functions_0|redist3|delay_signals[0][16] .power_up = "low";

dffeas \fp_functions_0|redist3|delay_signals[0][17] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][17]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist3|delay_signals[0][17]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist3|delay_signals[0][17] .is_wysiwyg = "true";
defparam \fp_functions_0|redist3|delay_signals[0][17] .power_up = "low";

dffeas \fp_functions_0|redist3|delay_signals[0][18] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][18]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist3|delay_signals[0][18]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist3|delay_signals[0][18] .is_wysiwyg = "true";
defparam \fp_functions_0|redist3|delay_signals[0][18] .power_up = "low";

dffeas \fp_functions_0|redist3|delay_signals[0][20] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][20]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist3|delay_signals[0][20]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist3|delay_signals[0][20] .is_wysiwyg = "true";
defparam \fp_functions_0|redist3|delay_signals[0][20] .power_up = "low";

dffeas \fp_functions_0|redist3|delay_signals[0][21] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][21]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist3|delay_signals[0][21]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist3|delay_signals[0][21] .is_wysiwyg = "true";
defparam \fp_functions_0|redist3|delay_signals[0][21] .power_up = "low";

dffeas \fp_functions_0|redist3|delay_signals[0][22] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][22]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist3|delay_signals[0][22]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist3|delay_signals[0][22] .is_wysiwyg = "true";
defparam \fp_functions_0|redist3|delay_signals[0][22] .power_up = "low";

dffeas \fp_functions_0|redist3|delay_signals[0][23] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][23]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist3|delay_signals[0][23]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist3|delay_signals[0][23] .is_wysiwyg = "true";
defparam \fp_functions_0|redist3|delay_signals[0][23] .power_up = "low";

dffeas \fp_functions_0|redist3|delay_signals[0][24] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][24]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist3|delay_signals[0][24]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist3|delay_signals[0][24] .is_wysiwyg = "true";
defparam \fp_functions_0|redist3|delay_signals[0][24] .power_up = "low";

dffeas \fp_functions_0|redist3|delay_signals[0][7] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][7]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist3|delay_signals[0][7]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist3|delay_signals[0][7] .is_wysiwyg = "true";
defparam \fp_functions_0|redist3|delay_signals[0][7] .power_up = "low";

dffeas \fp_functions_0|redist3|delay_signals[0][12] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][12]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist3|delay_signals[0][12]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist3|delay_signals[0][12] .is_wysiwyg = "true";
defparam \fp_functions_0|redist3|delay_signals[0][12] .power_up = "low";

dffeas \fp_functions_0|redist3|delay_signals[0][13] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][13]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist3|delay_signals[0][13]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist3|delay_signals[0][13] .is_wysiwyg = "true";
defparam \fp_functions_0|redist3|delay_signals[0][13] .power_up = "low";

dffeas \fp_functions_0|redist3|delay_signals[0][8] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][8]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist3|delay_signals[0][8]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist3|delay_signals[0][8] .is_wysiwyg = "true";
defparam \fp_functions_0|redist3|delay_signals[0][8] .power_up = "low";

dffeas \fp_functions_0|redist3|delay_signals[0][9] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][9]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist3|delay_signals[0][9]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist3|delay_signals[0][9] .is_wysiwyg = "true";
defparam \fp_functions_0|redist3|delay_signals[0][9] .power_up = "low";

dffeas \fp_functions_0|redist3|delay_signals[0][10] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][10]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist3|delay_signals[0][10]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist3|delay_signals[0][10] .is_wysiwyg = "true";
defparam \fp_functions_0|redist3|delay_signals[0][10] .power_up = "low";

dffeas \fp_functions_0|redist3|delay_signals[0][11] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][11]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist3|delay_signals[0][11]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist3|delay_signals[0][11] .is_wysiwyg = "true";
defparam \fp_functions_0|redist3|delay_signals[0][11] .power_up = "low";

dffeas \fp_functions_0|redist3|delay_signals[0][2] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][2]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist3|delay_signals[0][2]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist3|delay_signals[0][2] .is_wysiwyg = "true";
defparam \fp_functions_0|redist3|delay_signals[0][2] .power_up = "low";

dffeas \fp_functions_0|redist3|delay_signals[0][3] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][3]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist3|delay_signals[0][3]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist3|delay_signals[0][3] .is_wysiwyg = "true";
defparam \fp_functions_0|redist3|delay_signals[0][3] .power_up = "low";

dffeas \fp_functions_0|redist3|delay_signals[0][4] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][4]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist3|delay_signals[0][4]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist3|delay_signals[0][4] .is_wysiwyg = "true";
defparam \fp_functions_0|redist3|delay_signals[0][4] .power_up = "low";

dffeas \fp_functions_0|redist3|delay_signals[0][5] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][5]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist3|delay_signals[0][5]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist3|delay_signals[0][5] .is_wysiwyg = "true";
defparam \fp_functions_0|redist3|delay_signals[0][5] .power_up = "low";

dffeas \fp_functions_0|redist3|delay_signals[0][6] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][6]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist3|delay_signals[0][6]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist3|delay_signals[0][6] .is_wysiwyg = "true";
defparam \fp_functions_0|redist3|delay_signals[0][6] .power_up = "low";

dffeas \fp_functions_0|redist18|delay_signals[6][0] (
	.clk(clk),
	.d(\fp_functions_0|redist18|delay_signals[7][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist18|delay_signals[6][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist18|delay_signals[6][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist18|delay_signals[6][0] .power_up = "low";

dffeas \fp_functions_0|redist17|delay_signals[6][0] (
	.clk(clk),
	.d(\fp_functions_0|redist17|delay_signals[7][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist17|delay_signals[6][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist17|delay_signals[6][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist17|delay_signals[6][0] .power_up = "low";

dffeas \fp_functions_0|redist20|delay_signals[6][0] (
	.clk(clk),
	.d(\fp_functions_0|redist20|delay_signals[7][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist20|delay_signals[6][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist20|delay_signals[6][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist20|delay_signals[6][0] .power_up = "low";

dffeas \fp_functions_0|redist21|delay_signals[6][0] (
	.clk(clk),
	.d(\fp_functions_0|redist21|delay_signals[7][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist21|delay_signals[6][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist21|delay_signals[6][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist21|delay_signals[6][0] .power_up = "low";

dffeas \fp_functions_0|redist16|delay_signals[6][0] (
	.clk(clk),
	.d(\fp_functions_0|redist16|delay_signals[7][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist16|delay_signals[6][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist16|delay_signals[6][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist16|delay_signals[6][0] .power_up = "low";

dffeas \fp_functions_0|redist19|delay_signals[6][0] (
	.clk(clk),
	.d(\fp_functions_0|redist19|delay_signals[7][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist19|delay_signals[6][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist19|delay_signals[6][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist19|delay_signals[6][0] .power_up = "low";

dffeas \fp_functions_0|redist11|delay_signals[0][64] (
	.clk(clk),
	.d(\fp_functions_0|add_5~49_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist11|delay_signals[0][64]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist11|delay_signals[0][64] .is_wysiwyg = "true";
defparam \fp_functions_0|redist11|delay_signals[0][64] .power_up = "low";

dffeas \fp_functions_0|redist0|delay_signals[0][29] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][29]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist0|delay_signals[0][29]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist0|delay_signals[0][29] .is_wysiwyg = "true";
defparam \fp_functions_0|redist0|delay_signals[0][29] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][29] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][2]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][29]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][29] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][29] .power_up = "low";

dffeas \fp_functions_0|redist0|delay_signals[0][30] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][30]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist0|delay_signals[0][30]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist0|delay_signals[0][30] .is_wysiwyg = "true";
defparam \fp_functions_0|redist0|delay_signals[0][30] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][30] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][3]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][30]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][30] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][30] .power_up = "low";

dffeas \fp_functions_0|redist0|delay_signals[0][31] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][31]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist0|delay_signals[0][31]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist0|delay_signals[0][31] .is_wysiwyg = "true";
defparam \fp_functions_0|redist0|delay_signals[0][31] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][31] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][4]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][31]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][31] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][31] .power_up = "low";

dffeas \fp_functions_0|redist0|delay_signals[0][32] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][32]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist0|delay_signals[0][32]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist0|delay_signals[0][32] .is_wysiwyg = "true";
defparam \fp_functions_0|redist0|delay_signals[0][32] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][32] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][5]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][32]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][32] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][32] .power_up = "low";

dffeas \fp_functions_0|redist0|delay_signals[0][33] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][33]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist0|delay_signals[0][33]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist0|delay_signals[0][33] .is_wysiwyg = "true";
defparam \fp_functions_0|redist0|delay_signals[0][33] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][33] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][6]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][33]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][33] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][33] .power_up = "low";

dffeas \fp_functions_0|redist0|delay_signals[0][34] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][34]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist0|delay_signals[0][34]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist0|delay_signals[0][34] .is_wysiwyg = "true";
defparam \fp_functions_0|redist0|delay_signals[0][34] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][34] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][7]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][34]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][34] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][34] .power_up = "low";

dffeas \fp_functions_0|redist0|delay_signals[0][35] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][35]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist0|delay_signals[0][35]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist0|delay_signals[0][35] .is_wysiwyg = "true";
defparam \fp_functions_0|redist0|delay_signals[0][35] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][35] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][8]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][35]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][35] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][35] .power_up = "low";

dffeas \fp_functions_0|redist0|delay_signals[0][36] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][36]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist0|delay_signals[0][36]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist0|delay_signals[0][36] .is_wysiwyg = "true";
defparam \fp_functions_0|redist0|delay_signals[0][36] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][36] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][9]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][36]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][36] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][36] .power_up = "low";

dffeas \fp_functions_0|redist0|delay_signals[0][37] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][37]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist0|delay_signals[0][37]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist0|delay_signals[0][37] .is_wysiwyg = "true";
defparam \fp_functions_0|redist0|delay_signals[0][37] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][37] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][10]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][37]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][37] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][37] .power_up = "low";

dffeas \fp_functions_0|redist0|delay_signals[0][38] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][38]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist0|delay_signals[0][38]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist0|delay_signals[0][38] .is_wysiwyg = "true";
defparam \fp_functions_0|redist0|delay_signals[0][38] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][38] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][11]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][38]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][38] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][38] .power_up = "low";

dffeas \fp_functions_0|redist0|delay_signals[0][39] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][39]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist0|delay_signals[0][39]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist0|delay_signals[0][39] .is_wysiwyg = "true";
defparam \fp_functions_0|redist0|delay_signals[0][39] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][39] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][12]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][39]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][39] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][39] .power_up = "low";

dffeas \fp_functions_0|redist0|delay_signals[0][40] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][40]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist0|delay_signals[0][40]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist0|delay_signals[0][40] .is_wysiwyg = "true";
defparam \fp_functions_0|redist0|delay_signals[0][40] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][40] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][13]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][40]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][40] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][40] .power_up = "low";

dffeas \fp_functions_0|redist0|delay_signals[0][41] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][41]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist0|delay_signals[0][41]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist0|delay_signals[0][41] .is_wysiwyg = "true";
defparam \fp_functions_0|redist0|delay_signals[0][41] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][41] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][14]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][41]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][41] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][41] .power_up = "low";

dffeas \fp_functions_0|redist0|delay_signals[0][42] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][42]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist0|delay_signals[0][42]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist0|delay_signals[0][42] .is_wysiwyg = "true";
defparam \fp_functions_0|redist0|delay_signals[0][42] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][42] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][15]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][42]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][42] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][42] .power_up = "low";

dffeas \fp_functions_0|redist0|delay_signals[0][43] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][43]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist0|delay_signals[0][43]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist0|delay_signals[0][43] .is_wysiwyg = "true";
defparam \fp_functions_0|redist0|delay_signals[0][43] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][43] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][16]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][43]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][43] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][43] .power_up = "low";

dffeas \fp_functions_0|redist0|delay_signals[0][44] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][44]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist0|delay_signals[0][44]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist0|delay_signals[0][44] .is_wysiwyg = "true";
defparam \fp_functions_0|redist0|delay_signals[0][44] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][44] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][17]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][44]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][44] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][44] .power_up = "low";

dffeas \fp_functions_0|redist0|delay_signals[0][45] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][45]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist0|delay_signals[0][45]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist0|delay_signals[0][45] .is_wysiwyg = "true";
defparam \fp_functions_0|redist0|delay_signals[0][45] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][45] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][18]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][45]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][45] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][45] .power_up = "low";

dffeas \fp_functions_0|redist0|delay_signals[0][46] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][46]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist0|delay_signals[0][46]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist0|delay_signals[0][46] .is_wysiwyg = "true";
defparam \fp_functions_0|redist0|delay_signals[0][46] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][46] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][19]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][46]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][46] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][46] .power_up = "low";

dffeas \fp_functions_0|redist0|delay_signals[0][47] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][47]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist0|delay_signals[0][47]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist0|delay_signals[0][47] .is_wysiwyg = "true";
defparam \fp_functions_0|redist0|delay_signals[0][47] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][47] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][20]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][47]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][47] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][47] .power_up = "low";

dffeas \fp_functions_0|redist0|delay_signals[0][48] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][48]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist0|delay_signals[0][48]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist0|delay_signals[0][48] .is_wysiwyg = "true";
defparam \fp_functions_0|redist0|delay_signals[0][48] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][48] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][21]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][48]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][48] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][48] .power_up = "low";

dffeas \fp_functions_0|redist0|delay_signals[0][49] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][49]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist0|delay_signals[0][49]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist0|delay_signals[0][49] .is_wysiwyg = "true";
defparam \fp_functions_0|redist0|delay_signals[0][49] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][49] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][22]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][49]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][49] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][49] .power_up = "low";

dffeas \fp_functions_0|redist0|delay_signals[0][50] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][50]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist0|delay_signals[0][50]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist0|delay_signals[0][50] .is_wysiwyg = "true";
defparam \fp_functions_0|redist0|delay_signals[0][50] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][50] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][23]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][50]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][50] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][50] .power_up = "low";

dffeas \fp_functions_0|redist0|delay_signals[0][51] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][51]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist0|delay_signals[0][51]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist0|delay_signals[0][51] .is_wysiwyg = "true";
defparam \fp_functions_0|redist0|delay_signals[0][51] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][51] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][24]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][51]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][51] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][51] .power_up = "low";

dffeas \fp_functions_0|redist0|delay_signals[0][52] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][52]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist0|delay_signals[0][52]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist0|delay_signals[0][52] .is_wysiwyg = "true";
defparam \fp_functions_0|redist0|delay_signals[0][52] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][52] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][25]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][52]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][52] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][52] .power_up = "low";

dffeas \fp_functions_0|redist0|delay_signals[0][53] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][53]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist0|delay_signals[0][53]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist0|delay_signals[0][53] .is_wysiwyg = "true";
defparam \fp_functions_0|redist0|delay_signals[0][53] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][53] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][26]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][53]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][53] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][53] .power_up = "low";

dffeas \fp_functions_0|redist0|delay_signals[0][54] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][54]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist0|delay_signals[0][54]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist0|delay_signals[0][54] .is_wysiwyg = "true";
defparam \fp_functions_0|redist0|delay_signals[0][54] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][54] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][27]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][54]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][54] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][54] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][55] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][28]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][55]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][55] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][55] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][56] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][29]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][56]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][56] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][56] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][57] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][30]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][57]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][57] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][57] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][58] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][31]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][58]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][58] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][58] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][59] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][32]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][59]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][59] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][59] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][60] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][33]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][60]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][60] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][60] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][61] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][34]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][61]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][61] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][61] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][62] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][35]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][62]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][62] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][62] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][63] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][36]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][63]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][63] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][63] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][64] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][37]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][64]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][64] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][64] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][65] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][38]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][65]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][65] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][65] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][66] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][39]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][66]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][66] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][66] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][67] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][40]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][67]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][67] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][67] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][68] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][41]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][68]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][68] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][68] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][69] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][42]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][69]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][69] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][69] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][70] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][43]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][70]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][70] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][70] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][71] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][44]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][71]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][71] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][71] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][72] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][45]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][72]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][72] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][72] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][73] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][46]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][73]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][73] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][73] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][74] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][47]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][74]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][74] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][74] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][75] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][48]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][75]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][75] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][75] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][76] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][49]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][76]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][76] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][76] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][77] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][50]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][77]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][77] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][77] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][78] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][51]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][78]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][78] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][78] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][79] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][52]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][79]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][79] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][79] .power_up = "low";

dffeas \fp_functions_0|redist15_wraddr_q[0] (
	.clk(clk),
	.d(\fp_functions_0|i5779~0_combout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\fp_functions_0|redist15_wraddr_q[0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist15_wraddr_q[0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist15_wraddr_q[0] .power_up = "low";

dffeas \fp_functions_0|redist15_wraddr_q[1] (
	.clk(clk),
	.d(\fp_functions_0|i5779~1_combout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\fp_functions_0|redist15_wraddr_q[1]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist15_wraddr_q[1] .is_wysiwyg = "true";
defparam \fp_functions_0|redist15_wraddr_q[1] .power_up = "low";

dffeas \fp_functions_0|redist15_inputreg|delay_signals[0][0] (
	.clk(clk),
	.d(\fp_functions_0|expSum_uid44_fpMulTest_o[0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist15_inputreg|delay_signals[0][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist15_inputreg|delay_signals[0][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist15_inputreg|delay_signals[0][0] .power_up = "low";

dffeas \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|rdaddr_reg[0] (
	.clk(clk),
	.d(\fp_functions_0|i5779~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|rdaddr_reg[0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|rdaddr_reg[0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|rdaddr_reg[0] .power_up = "low";

dffeas \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|rdaddr_reg[1] (
	.clk(clk),
	.d(\fp_functions_0|i5779~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|rdaddr_reg[1]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|rdaddr_reg[1] .is_wysiwyg = "true";
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|rdaddr_reg[1] .power_up = "low";

dffeas \fp_functions_0|redist15_cmpReg_q[0] (
	.clk(clk),
	.d(\fp_functions_0|reduce_nor_8~combout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist15_cmpReg_q[0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist15_cmpReg_q[0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist15_cmpReg_q[0] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|redist15_sticky_ena_q[0]~0 (
	.dataa(!en[0]),
	.datab(!\fp_functions_0|redist15_sticky_ena_q[0]~q ),
	.datac(!\fp_functions_0|redist15_cmpReg_q[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|redist15_sticky_ena_q[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|redist15_sticky_ena_q[0]~0 .extended_lut = "off";
defparam \fp_functions_0|redist15_sticky_ena_q[0]~0 .lut_mask = 64'h3737373737373737;
defparam \fp_functions_0|redist15_sticky_ena_q[0]~0 .shared_arith = "off";

dffeas \fp_functions_0|redist14|delay_signals[7][0] (
	.clk(clk),
	.d(\fp_functions_0|redist14|delay_signals[8][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist14|delay_signals[7][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist14|delay_signals[7][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist14|delay_signals[7][0] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][27] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][27] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][27]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][27] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][27] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][0] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][0] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][0] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][0] .power_up = "low";

dffeas \fp_functions_0|redist0|delay_signals[0][26] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][26]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist0|delay_signals[0][26]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist0|delay_signals[0][26] .is_wysiwyg = "true";
defparam \fp_functions_0|redist0|delay_signals[0][26] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][26] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][53]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][26]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][26] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][26] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][28] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][28] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][28]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][28] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][28] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][1] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][1] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][1]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][1] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][1] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][53] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][53] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][53]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][53] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][53] .power_up = "low";

dffeas \fp_functions_0|redist0|delay_signals[0][23] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][23]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist0|delay_signals[0][23]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist0|delay_signals[0][23] .is_wysiwyg = "true";
defparam \fp_functions_0|redist0|delay_signals[0][23] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][23] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][50]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][23]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][23] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][23] .power_up = "low";

dffeas \fp_functions_0|redist0|delay_signals[0][24] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][24]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist0|delay_signals[0][24]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist0|delay_signals[0][24] .is_wysiwyg = "true";
defparam \fp_functions_0|redist0|delay_signals[0][24] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][24] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][51]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][24]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][24] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][24] .power_up = "low";

dffeas \fp_functions_0|redist0|delay_signals[0][25] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][25]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist0|delay_signals[0][25]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist0|delay_signals[0][25] .is_wysiwyg = "true";
defparam \fp_functions_0|redist0|delay_signals[0][25] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][25] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][52]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][25]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][25] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][25] .power_up = "low";

dffeas \fp_functions_0|redist0|delay_signals[0][16] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][16]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist0|delay_signals[0][16]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist0|delay_signals[0][16] .is_wysiwyg = "true";
defparam \fp_functions_0|redist0|delay_signals[0][16] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][16] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][43]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][16]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][16] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][16] .power_up = "low";

dffeas \fp_functions_0|redist0|delay_signals[0][21] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][21]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist0|delay_signals[0][21]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist0|delay_signals[0][21] .is_wysiwyg = "true";
defparam \fp_functions_0|redist0|delay_signals[0][21] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][21] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][48]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][21]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][21] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][21] .power_up = "low";

dffeas \fp_functions_0|redist0|delay_signals[0][22] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][22]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist0|delay_signals[0][22]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist0|delay_signals[0][22] .is_wysiwyg = "true";
defparam \fp_functions_0|redist0|delay_signals[0][22] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][22] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][49]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][22]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][22] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][22] .power_up = "low";

dffeas \fp_functions_0|redist0|delay_signals[0][17] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][17]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist0|delay_signals[0][17]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist0|delay_signals[0][17] .is_wysiwyg = "true";
defparam \fp_functions_0|redist0|delay_signals[0][17] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][17] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][44]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][17]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][17] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][17] .power_up = "low";

dffeas \fp_functions_0|redist0|delay_signals[0][18] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][18]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist0|delay_signals[0][18]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist0|delay_signals[0][18] .is_wysiwyg = "true";
defparam \fp_functions_0|redist0|delay_signals[0][18] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][18] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][45]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][18]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][18] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][18] .power_up = "low";

dffeas \fp_functions_0|redist0|delay_signals[0][19] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][19]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist0|delay_signals[0][19]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist0|delay_signals[0][19] .is_wysiwyg = "true";
defparam \fp_functions_0|redist0|delay_signals[0][19] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][19] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][46]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][19]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][19] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][19] .power_up = "low";

dffeas \fp_functions_0|redist0|delay_signals[0][20] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][20]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist0|delay_signals[0][20]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist0|delay_signals[0][20] .is_wysiwyg = "true";
defparam \fp_functions_0|redist0|delay_signals[0][20] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][20] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][47]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][20]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][20] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][20] .power_up = "low";

dffeas \fp_functions_0|redist0|delay_signals[0][11] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][11]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist0|delay_signals[0][11]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist0|delay_signals[0][11] .is_wysiwyg = "true";
defparam \fp_functions_0|redist0|delay_signals[0][11] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][11] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][38]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][11]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][11] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][11] .power_up = "low";

dffeas \fp_functions_0|redist0|delay_signals[0][12] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][12]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist0|delay_signals[0][12]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist0|delay_signals[0][12] .is_wysiwyg = "true";
defparam \fp_functions_0|redist0|delay_signals[0][12] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][12] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][39]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][12]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][12] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][12] .power_up = "low";

dffeas \fp_functions_0|redist0|delay_signals[0][13] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][13]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist0|delay_signals[0][13]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist0|delay_signals[0][13] .is_wysiwyg = "true";
defparam \fp_functions_0|redist0|delay_signals[0][13] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][13] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][40]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][13]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][13] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][13] .power_up = "low";

dffeas \fp_functions_0|redist0|delay_signals[0][14] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][14]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist0|delay_signals[0][14]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist0|delay_signals[0][14] .is_wysiwyg = "true";
defparam \fp_functions_0|redist0|delay_signals[0][14] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][14] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][41]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][14]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][14] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][14] .power_up = "low";

dffeas \fp_functions_0|redist0|delay_signals[0][15] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][15]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist0|delay_signals[0][15]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist0|delay_signals[0][15] .is_wysiwyg = "true";
defparam \fp_functions_0|redist0|delay_signals[0][15] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][15] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][42]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][15]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][15] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][15] .power_up = "low";

dffeas \fp_functions_0|redist0|delay_signals[0][4] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][4]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist0|delay_signals[0][4]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist0|delay_signals[0][4] .is_wysiwyg = "true";
defparam \fp_functions_0|redist0|delay_signals[0][4] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][4] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][31]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][4]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][4] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][4] .power_up = "low";

dffeas \fp_functions_0|redist0|delay_signals[0][10] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][10]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist0|delay_signals[0][10]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist0|delay_signals[0][10] .is_wysiwyg = "true";
defparam \fp_functions_0|redist0|delay_signals[0][10] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][10] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][37]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][10]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][10] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][10] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][26] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][26] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][26]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][26] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][26] .power_up = "low";

dffeas \fp_functions_0|redist0|delay_signals[0][0] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist0|delay_signals[0][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist0|delay_signals[0][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist0|delay_signals[0][0] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][0] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][27]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][0] .power_up = "low";

dffeas \fp_functions_0|redist0|delay_signals[0][1] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][1]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist0|delay_signals[0][1]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist0|delay_signals[0][1] .is_wysiwyg = "true";
defparam \fp_functions_0|redist0|delay_signals[0][1] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][1] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][28]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][1]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][1] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][1] .power_up = "low";

dffeas \fp_functions_0|redist0|delay_signals[0][2] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][2]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist0|delay_signals[0][2]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist0|delay_signals[0][2] .is_wysiwyg = "true";
defparam \fp_functions_0|redist0|delay_signals[0][2] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][2] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][29]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][2]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][2] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][2] .power_up = "low";

dffeas \fp_functions_0|redist0|delay_signals[0][3] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][3]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist0|delay_signals[0][3]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist0|delay_signals[0][3] .is_wysiwyg = "true";
defparam \fp_functions_0|redist0|delay_signals[0][3] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][3] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][30]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][3]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][3] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][3] .power_up = "low";

dffeas \fp_functions_0|redist0|delay_signals[0][5] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][5]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist0|delay_signals[0][5]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist0|delay_signals[0][5] .is_wysiwyg = "true";
defparam \fp_functions_0|redist0|delay_signals[0][5] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][5] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][32]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][5]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][5] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][5] .power_up = "low";

dffeas \fp_functions_0|redist0|delay_signals[0][6] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][6]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist0|delay_signals[0][6]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist0|delay_signals[0][6] .is_wysiwyg = "true";
defparam \fp_functions_0|redist0|delay_signals[0][6] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][6] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][33]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][6]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][6] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][6] .power_up = "low";

dffeas \fp_functions_0|redist0|delay_signals[0][7] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][7]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist0|delay_signals[0][7]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist0|delay_signals[0][7] .is_wysiwyg = "true";
defparam \fp_functions_0|redist0|delay_signals[0][7] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][7] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][34]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][7]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][7] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][7] .power_up = "low";

dffeas \fp_functions_0|redist0|delay_signals[0][8] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][8]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist0|delay_signals[0][8]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist0|delay_signals[0][8] .is_wysiwyg = "true";
defparam \fp_functions_0|redist0|delay_signals[0][8] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][8] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][35]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][8]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][8] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][8] .power_up = "low";

dffeas \fp_functions_0|redist0|delay_signals[0][9] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][9]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist0|delay_signals[0][9]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist0|delay_signals[0][9] .is_wysiwyg = "true";
defparam \fp_functions_0|redist0|delay_signals[0][9] .power_up = "low";

dffeas \fp_functions_0|redist2|delay_signals[0][9] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][36]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist2|delay_signals[0][9]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist2|delay_signals[0][9] .is_wysiwyg = "true";
defparam \fp_functions_0|redist2|delay_signals[0][9] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][19] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][19] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][19]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][19] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][19] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][25] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][25] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][25]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][25] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][25] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][14] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][14] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][14]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][14] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][14] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][15] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][15] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][15]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][15] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][15] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][16] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][16] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][16]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][16] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][16] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][17] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][17] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][17]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][17] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][17] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][18] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][18] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][18]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][18] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][18] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][20] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][20] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][20]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][20] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][20] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][21] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][21] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][21]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][21] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][21] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][22] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][22] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][22]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][22] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][22] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][23] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][23] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][23]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][23] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][23] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][24] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][24] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][24]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][24] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][24] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][7] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][7] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][7]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][7] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][7] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][12] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][12] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][12]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][12] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][12] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][13] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][13] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][13]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][13] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][13] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][8] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][8] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][8]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][8] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][8] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][9] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][9] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][9]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][9] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][9] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][10] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][10] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][10]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][10] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][10] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][11] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][11] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][11]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][11] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][11] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][2] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][2] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][2]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][2] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][2] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][3] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][3] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][3]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][3] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][3] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][4] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][4] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][4]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][4] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][4] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][5] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][5] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][5]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][5] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][5] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][6] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][6] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][6]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][6] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][6] .power_up = "low";

dffeas \fp_functions_0|redist18|delay_signals[7][0] (
	.clk(clk),
	.d(\fp_functions_0|excZ_y_uid29_fpMulTest_delay|delay_signals[0][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist18|delay_signals[7][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist18|delay_signals[7][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist18|delay_signals[7][0] .power_up = "low";

dffeas \fp_functions_0|redist17|delay_signals[7][0] (
	.clk(clk),
	.d(\fp_functions_0|expXIsMax_uid30_fpMulTest_delay|delay_signals[0][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist17|delay_signals[7][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist17|delay_signals[7][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist17|delay_signals[7][0] .power_up = "low";

dffeas \fp_functions_0|redist20|delay_signals[7][0] (
	.clk(clk),
	.d(\fp_functions_0|expXIsMax_uid16_fpMulTest_delay|delay_signals[0][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist20|delay_signals[7][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist20|delay_signals[7][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist20|delay_signals[7][0] .power_up = "low";

dffeas \fp_functions_0|redist21|delay_signals[7][0] (
	.clk(clk),
	.d(\fp_functions_0|excZ_x_uid15_fpMulTest_delay|delay_signals[0][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist21|delay_signals[7][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist21|delay_signals[7][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist21|delay_signals[7][0] .power_up = "low";

dffeas \fp_functions_0|redist16|delay_signals[7][0] (
	.clk(clk),
	.d(\fp_functions_0|fracXIsZero_uid31_fpMulTest_delay|delay_signals[0][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist16|delay_signals[7][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist16|delay_signals[7][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist16|delay_signals[7][0] .power_up = "low";

dffeas \fp_functions_0|redist19|delay_signals[7][0] (
	.clk(clk),
	.d(\fp_functions_0|fracXIsZero_uid17_fpMulTest_delay|delay_signals[0][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist19|delay_signals[7][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist19|delay_signals[7][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist19|delay_signals[7][0] .power_up = "low";

dffeas \fp_functions_0|redist15_outputreg|delay_signals[0][11] (
	.clk(clk),
	.d(\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[11]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist15_outputreg|delay_signals[0][11]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist15_outputreg|delay_signals[0][11] .is_wysiwyg = "true";
defparam \fp_functions_0|redist15_outputreg|delay_signals[0][11] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][29] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][29] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][29]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][29] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][29] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][2] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][2] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][2]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][2] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][2] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][30] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][30] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][30]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][30] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][30] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][3] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][3] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][3]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][3] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][3] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][31] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][31] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][31]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][31] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][31] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][4] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][4] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][4]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][4] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][4] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][32] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][32] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][32]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][32] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][32] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][5] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][5] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][5]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][5] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][5] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][33] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][33] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][33]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][33] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][33] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][6] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][6] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][6]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][6] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][6] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][34] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][34] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][34]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][34] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][34] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][7] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][7] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][7]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][7] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][7] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][35] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][35] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][35]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][35] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][35] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][8] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][8] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][8]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][8] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][8] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][36] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][36] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][36]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][36] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][36] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][9] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][9] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][9]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][9] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][9] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][37] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][37] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][37]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][37] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][37] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][10] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][10] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][10]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][10] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][10] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][38] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][38] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][38]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][38] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][38] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][11] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][11] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][11]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][11] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][11] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][39] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][39] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][39]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][39] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][39] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][12] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][12] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][12]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][12] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][12] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][40] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][40] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][40]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][40] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][40] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][13] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][13] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][13]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][13] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][13] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][41] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][41] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][41]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][41] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][41] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][14] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][14] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][14]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][14] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][14] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][42] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][42] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][42]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][42] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][42] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][15] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][15] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][15]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][15] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][15] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][43] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][43] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][43]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][43] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][43] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][16] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][16] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][16]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][16] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][16] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][44] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][44] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][44]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][44] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][44] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][17] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][17] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][17]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][17] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][17] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][45] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][45] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][45]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][45] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][45] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][18] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][18] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][18]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][18] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][18] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][46] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][46] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][46]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][46] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][46] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][19] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][19] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][19]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][19] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][19] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][47] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][47] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][47]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][47] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][47] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][20] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][20] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][20]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][20] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][20] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][48] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][48] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][48]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][48] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][48] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][21] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][21] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][21]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][21] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][21] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][49] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][49] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][49]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][49] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][49] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][22] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][22] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][22]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][22] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][22] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][50] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][50] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][50]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][50] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][50] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][23] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][23] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][23]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][23] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][23] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][51] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][51] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][51]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][51] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][51] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][24] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][24] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][24]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][24] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][24] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][52] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][52] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][52]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][52] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][52] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][25] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][25] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][25]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][25] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][25] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][53] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][53] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][53]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][53] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][53] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][26] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][26] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][26]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][26] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][26] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][54] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][54] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][54]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][54] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][54] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][27] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][27] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][27]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][27] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][27] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][28] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][28] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][28]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][28] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][28] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][29] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][29] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][29]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][29] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][29] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][30] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][30] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][30]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][30] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][30] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][31] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][31] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][31]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][31] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][31] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][32] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][32] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][32]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][32] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][32] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][33] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][33] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][33]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][33] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][33] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][34] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][34] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][34]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][34] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][34] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][35] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][35] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][35]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][35] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][35] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][36] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][36] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][36]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][36] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][36] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][37] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][37] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][37]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][37] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][37] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][38] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][38] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][38]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][38] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][38] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][39] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][39] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][39]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][39] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][39] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][40] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][40] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][40]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][40] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][40] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][41] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][41] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][41]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][41] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][41] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][42] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][42] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][42]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][42] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][42] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][43] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][43] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][43]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][43] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][43] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][44] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][44] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][44]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][44] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][44] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][45] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][45] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][45]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][45] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][45] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][46] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][46] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][46]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][46] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][46] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][47] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][47] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][47]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][47] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][47] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][48] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][48] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][48]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][48] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][48] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][49] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][49] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][49]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][49] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][49] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][50] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][50] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][50]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][50] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][50] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][51] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][51] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][51]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][51] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][51] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][52] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_y[0][52] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][52]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][52] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_s[0][52] .power_up = "low";

dffeas \fp_functions_0|redist15_rdcnt_i[0] (
	.clk(clk),
	.d(\fp_functions_0|redist15_rdcnt_i[0]~0_combout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\fp_functions_0|redist15_rdcnt_i[0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist15_rdcnt_i[0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist15_rdcnt_i[0] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|i5779~0 (
	.dataa(!en[0]),
	.datab(!\fp_functions_0|redist15_wraddr_q[0]~q ),
	.datac(!\fp_functions_0|redist15_rdcnt_i[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|i5779~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|i5779~0 .extended_lut = "off";
defparam \fp_functions_0|i5779~0 .lut_mask = 64'h7272727272727272;
defparam \fp_functions_0|i5779~0 .shared_arith = "off";

dffeas \fp_functions_0|redist15_rdcnt_i[1] (
	.clk(clk),
	.d(\fp_functions_0|i5766~0_combout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist15_rdcnt_i[1]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist15_rdcnt_i[1] .is_wysiwyg = "true";
defparam \fp_functions_0|redist15_rdcnt_i[1] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|i5779~1 (
	.dataa(!en[0]),
	.datab(!\fp_functions_0|redist15_wraddr_q[1]~q ),
	.datac(!\fp_functions_0|redist15_rdcnt_i[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|i5779~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|i5779~1 .extended_lut = "off";
defparam \fp_functions_0|i5779~1 .lut_mask = 64'h2727272727272727;
defparam \fp_functions_0|i5779~1 .shared_arith = "off";

dffeas \fp_functions_0|expSum_uid44_fpMulTest_o[0] (
	.clk(clk),
	.d(\fp_functions_0|add_4~1_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|expSum_uid44_fpMulTest_o[0]~q ),
	.prn(vcc));
defparam \fp_functions_0|expSum_uid44_fpMulTest_o[0] .is_wysiwyg = "true";
defparam \fp_functions_0|expSum_uid44_fpMulTest_o[0] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|reduce_nor_8 (
	.dataa(!en[0]),
	.datab(!\fp_functions_0|redist15_wraddr_q[0]~q ),
	.datac(!\fp_functions_0|redist15_wraddr_q[1]~q ),
	.datad(!\fp_functions_0|redist15_rdcnt_i[0]~q ),
	.datae(!\fp_functions_0|redist15_rdcnt_i[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|reduce_nor_8~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|reduce_nor_8 .extended_lut = "off";
defparam \fp_functions_0|reduce_nor_8 .lut_mask = 64'h0808085D0808085D;
defparam \fp_functions_0|reduce_nor_8 .shared_arith = "off";

dffeas \fp_functions_0|redist15_inputreg|delay_signals[0][1] (
	.clk(clk),
	.d(\fp_functions_0|expSum_uid44_fpMulTest_o[1]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist15_inputreg|delay_signals[0][1]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist15_inputreg|delay_signals[0][1] .is_wysiwyg = "true";
defparam \fp_functions_0|redist15_inputreg|delay_signals[0][1] .power_up = "low";

dffeas \fp_functions_0|redist15_inputreg|delay_signals[0][2] (
	.clk(clk),
	.d(\fp_functions_0|expSum_uid44_fpMulTest_o[2]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist15_inputreg|delay_signals[0][2]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist15_inputreg|delay_signals[0][2] .is_wysiwyg = "true";
defparam \fp_functions_0|redist15_inputreg|delay_signals[0][2] .power_up = "low";

dffeas \fp_functions_0|redist15_inputreg|delay_signals[0][3] (
	.clk(clk),
	.d(\fp_functions_0|expSum_uid44_fpMulTest_o[3]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist15_inputreg|delay_signals[0][3]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist15_inputreg|delay_signals[0][3] .is_wysiwyg = "true";
defparam \fp_functions_0|redist15_inputreg|delay_signals[0][3] .power_up = "low";

dffeas \fp_functions_0|redist15_inputreg|delay_signals[0][4] (
	.clk(clk),
	.d(\fp_functions_0|expSum_uid44_fpMulTest_o[4]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist15_inputreg|delay_signals[0][4]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist15_inputreg|delay_signals[0][4] .is_wysiwyg = "true";
defparam \fp_functions_0|redist15_inputreg|delay_signals[0][4] .power_up = "low";

dffeas \fp_functions_0|redist15_inputreg|delay_signals[0][5] (
	.clk(clk),
	.d(\fp_functions_0|expSum_uid44_fpMulTest_o[5]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist15_inputreg|delay_signals[0][5]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist15_inputreg|delay_signals[0][5] .is_wysiwyg = "true";
defparam \fp_functions_0|redist15_inputreg|delay_signals[0][5] .power_up = "low";

dffeas \fp_functions_0|redist15_inputreg|delay_signals[0][6] (
	.clk(clk),
	.d(\fp_functions_0|expSum_uid44_fpMulTest_o[6]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist15_inputreg|delay_signals[0][6]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist15_inputreg|delay_signals[0][6] .is_wysiwyg = "true";
defparam \fp_functions_0|redist15_inputreg|delay_signals[0][6] .power_up = "low";

dffeas \fp_functions_0|redist15_inputreg|delay_signals[0][7] (
	.clk(clk),
	.d(\fp_functions_0|expSum_uid44_fpMulTest_o[7]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist15_inputreg|delay_signals[0][7]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist15_inputreg|delay_signals[0][7] .is_wysiwyg = "true";
defparam \fp_functions_0|redist15_inputreg|delay_signals[0][7] .power_up = "low";

dffeas \fp_functions_0|redist15_inputreg|delay_signals[0][8] (
	.clk(clk),
	.d(\fp_functions_0|expSum_uid44_fpMulTest_o[8]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist15_inputreg|delay_signals[0][8]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist15_inputreg|delay_signals[0][8] .is_wysiwyg = "true";
defparam \fp_functions_0|redist15_inputreg|delay_signals[0][8] .power_up = "low";

dffeas \fp_functions_0|redist15_inputreg|delay_signals[0][9] (
	.clk(clk),
	.d(\fp_functions_0|expSum_uid44_fpMulTest_o[9]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist15_inputreg|delay_signals[0][9]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist15_inputreg|delay_signals[0][9] .is_wysiwyg = "true";
defparam \fp_functions_0|redist15_inputreg|delay_signals[0][9] .power_up = "low";

dffeas \fp_functions_0|redist15_inputreg|delay_signals[0][10] (
	.clk(clk),
	.d(\fp_functions_0|expSum_uid44_fpMulTest_o[10]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist15_inputreg|delay_signals[0][10]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist15_inputreg|delay_signals[0][10] .is_wysiwyg = "true";
defparam \fp_functions_0|redist15_inputreg|delay_signals[0][10] .power_up = "low";

dffeas \fp_functions_0|redist14|delay_signals[8][0] (
	.clk(clk),
	.d(\fp_functions_0|signR_uid48_fpMulTest_delay|delay_signals[0][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist14|delay_signals[8][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist14|delay_signals[8][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist14|delay_signals[8][0] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][26] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][26] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][26]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][26] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][26] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][53] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][53] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][53]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][53] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][53] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][23] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][23] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][23]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][23] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][23] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][50] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][50] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][50]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][50] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][50] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][24] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][24] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][24]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][24] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][24] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][51] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][51] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][51]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][51] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][51] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][25] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][25] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][25]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][25] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][25] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][52] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][52] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][52]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][52] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][52] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][16] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][16] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][16]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][16] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][16] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][43] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][43] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][43]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][43] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][43] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][21] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][21] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][21]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][21] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][21] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][48] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][48] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][48]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][48] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][48] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][22] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][22] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][22]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][22] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][22] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][49] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][49] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][49]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][49] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][49] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][17] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][17] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][17]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][17] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][17] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][44] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][44] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][44]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][44] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][44] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][18] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][18] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][18]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][18] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][18] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][45] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][45] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][45]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][45] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][45] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][19] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][19] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][19]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][19] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][19] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][46] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][46] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][46]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][46] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][46] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][20] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][20] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][20]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][20] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][20] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][47] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][47] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][47]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][47] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][47] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][11] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][11] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][11]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][11] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][11] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][38] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][38] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][38]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][38] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][38] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][12] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][12] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][12]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][12] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][12] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][39] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][39] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][39]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][39] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][39] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][13] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][13] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][13]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][13] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][13] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][40] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][40] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][40]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][40] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][40] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][14] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][14] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][14]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][14] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][14] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][41] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][41] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][41]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][41] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][41] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][15] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][15] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][15]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][15] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][15] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][42] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][42] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][42]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][42] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][42] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][4] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][4] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][4]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][4] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][4] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][31] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][31] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][31]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][31] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][31] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][10] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][10] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][10]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][10] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][10] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][37] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][37] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][37]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][37] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][37] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][0] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][0] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][0] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][0] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][27] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][27] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][27]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][27] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][27] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][1] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][1] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][1]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][1] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][1] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][28] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][28] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][28]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][28] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][28] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][2] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][2] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][2]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][2] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][2] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][29] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][29] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][29]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][29] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][29] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][3] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][3] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][3]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][3] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][3] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][30] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][30] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][30]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][30] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][30] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][5] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][5] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][5]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][5] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][5] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][32] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][32] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][32]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][32] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][32] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][6] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][6] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][6]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][6] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][6] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][33] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][33] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][33]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][33] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][33] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][7] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][7] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][7]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][7] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][7] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][34] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][34] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][34]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][34] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][34] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][8] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][8] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][8]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][8] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][8] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][35] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][35] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][35]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][35] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][35] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][9] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_y[0][9] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][9]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][9] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_s[0][9] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][36] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_y[0][36] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][36]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][36] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_s[0][36] .power_up = "low";

dffeas \fp_functions_0|excZ_y_uid29_fpMulTest_delay|delay_signals[0][0] (
	.clk(clk),
	.d(\fp_functions_0|reduce_nor_2~combout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|excZ_y_uid29_fpMulTest_delay|delay_signals[0][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|excZ_y_uid29_fpMulTest_delay|delay_signals[0][0] .is_wysiwyg = "true";
defparam \fp_functions_0|excZ_y_uid29_fpMulTest_delay|delay_signals[0][0] .power_up = "low";

dffeas \fp_functions_0|expXIsMax_uid30_fpMulTest_delay|delay_signals[0][0] (
	.clk(clk),
	.d(\fp_functions_0|reduce_nor_4~combout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|expXIsMax_uid30_fpMulTest_delay|delay_signals[0][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|expXIsMax_uid30_fpMulTest_delay|delay_signals[0][0] .is_wysiwyg = "true";
defparam \fp_functions_0|expXIsMax_uid30_fpMulTest_delay|delay_signals[0][0] .power_up = "low";

dffeas \fp_functions_0|expXIsMax_uid16_fpMulTest_delay|delay_signals[0][0] (
	.clk(clk),
	.d(\fp_functions_0|reduce_nor_1~combout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|expXIsMax_uid16_fpMulTest_delay|delay_signals[0][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|expXIsMax_uid16_fpMulTest_delay|delay_signals[0][0] .is_wysiwyg = "true";
defparam \fp_functions_0|expXIsMax_uid16_fpMulTest_delay|delay_signals[0][0] .power_up = "low";

dffeas \fp_functions_0|excZ_x_uid15_fpMulTest_delay|delay_signals[0][0] (
	.clk(clk),
	.d(\fp_functions_0|reduce_nor_5~combout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|excZ_x_uid15_fpMulTest_delay|delay_signals[0][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|excZ_x_uid15_fpMulTest_delay|delay_signals[0][0] .is_wysiwyg = "true";
defparam \fp_functions_0|excZ_x_uid15_fpMulTest_delay|delay_signals[0][0] .power_up = "low";

dffeas \fp_functions_0|fracXIsZero_uid31_fpMulTest_delay|delay_signals[0][0] (
	.clk(clk),
	.d(\fp_functions_0|reduce_nor_3~combout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|fracXIsZero_uid31_fpMulTest_delay|delay_signals[0][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|fracXIsZero_uid31_fpMulTest_delay|delay_signals[0][0] .is_wysiwyg = "true";
defparam \fp_functions_0|fracXIsZero_uid31_fpMulTest_delay|delay_signals[0][0] .power_up = "low";

dffeas \fp_functions_0|fracXIsZero_uid17_fpMulTest_delay|delay_signals[0][0] (
	.clk(clk),
	.d(\fp_functions_0|reduce_nor_0~combout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|fracXIsZero_uid17_fpMulTest_delay|delay_signals[0][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|fracXIsZero_uid17_fpMulTest_delay|delay_signals[0][0] .is_wysiwyg = "true";
defparam \fp_functions_0|fracXIsZero_uid17_fpMulTest_delay|delay_signals[0][0] .power_up = "low";

dffeas \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[11] (
	.clk(clk),
	.d(\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_wire[11] ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\fp_functions_0|i5762~combout ),
	.q(\fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[11]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[11] .is_wysiwyg = "true";
defparam \fp_functions_0|redist15_mem_dmem|auto_generated|altsyncram1|dataout_reg[11] .power_up = "low";

dffeas \fp_functions_0|redist15_rdcnt_eq (
	.clk(clk),
	.d(\fp_functions_0|reduce_nor_9~combout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist15_rdcnt_eq~q ),
	.prn(vcc));
defparam \fp_functions_0|redist15_rdcnt_eq .is_wysiwyg = "true";
defparam \fp_functions_0|redist15_rdcnt_eq .power_up = "low";

twentynm_lcell_comb \fp_functions_0|redist15_rdcnt_i[0]~0 (
	.dataa(!en[0]),
	.datab(!\fp_functions_0|redist15_rdcnt_i[0]~q ),
	.datac(!\fp_functions_0|redist15_rdcnt_eq~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|redist15_rdcnt_i[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|redist15_rdcnt_i[0]~0 .extended_lut = "off";
defparam \fp_functions_0|redist15_rdcnt_i[0]~0 .lut_mask = 64'h6363636363636363;
defparam \fp_functions_0|redist15_rdcnt_i[0]~0 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|i5766~0 (
	.dataa(!\fp_functions_0|redist15_rdcnt_i[0]~q ),
	.datab(!\fp_functions_0|redist15_rdcnt_i[1]~q ),
	.datac(!\fp_functions_0|redist15_rdcnt_eq~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|i5766~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|i5766~0 .extended_lut = "off";
defparam \fp_functions_0|i5766~0 .lut_mask = 64'h9C9C9C9C9C9C9C9C;
defparam \fp_functions_0|i5766~0 .shared_arith = "off";

dffeas \fp_functions_0|expSum_uid44_fpMulTest_o[1] (
	.clk(clk),
	.d(\fp_functions_0|add_4~5_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|expSum_uid44_fpMulTest_o[1]~q ),
	.prn(vcc));
defparam \fp_functions_0|expSum_uid44_fpMulTest_o[1] .is_wysiwyg = "true";
defparam \fp_functions_0|expSum_uid44_fpMulTest_o[1] .power_up = "low";

dffeas \fp_functions_0|expSum_uid44_fpMulTest_o[2] (
	.clk(clk),
	.d(\fp_functions_0|add_4~9_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|expSum_uid44_fpMulTest_o[2]~q ),
	.prn(vcc));
defparam \fp_functions_0|expSum_uid44_fpMulTest_o[2] .is_wysiwyg = "true";
defparam \fp_functions_0|expSum_uid44_fpMulTest_o[2] .power_up = "low";

dffeas \fp_functions_0|expSum_uid44_fpMulTest_o[3] (
	.clk(clk),
	.d(\fp_functions_0|add_4~13_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|expSum_uid44_fpMulTest_o[3]~q ),
	.prn(vcc));
defparam \fp_functions_0|expSum_uid44_fpMulTest_o[3] .is_wysiwyg = "true";
defparam \fp_functions_0|expSum_uid44_fpMulTest_o[3] .power_up = "low";

dffeas \fp_functions_0|expSum_uid44_fpMulTest_o[4] (
	.clk(clk),
	.d(\fp_functions_0|add_4~17_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|expSum_uid44_fpMulTest_o[4]~q ),
	.prn(vcc));
defparam \fp_functions_0|expSum_uid44_fpMulTest_o[4] .is_wysiwyg = "true";
defparam \fp_functions_0|expSum_uid44_fpMulTest_o[4] .power_up = "low";

dffeas \fp_functions_0|expSum_uid44_fpMulTest_o[5] (
	.clk(clk),
	.d(\fp_functions_0|add_4~21_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|expSum_uid44_fpMulTest_o[5]~q ),
	.prn(vcc));
defparam \fp_functions_0|expSum_uid44_fpMulTest_o[5] .is_wysiwyg = "true";
defparam \fp_functions_0|expSum_uid44_fpMulTest_o[5] .power_up = "low";

dffeas \fp_functions_0|expSum_uid44_fpMulTest_o[6] (
	.clk(clk),
	.d(\fp_functions_0|add_4~25_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|expSum_uid44_fpMulTest_o[6]~q ),
	.prn(vcc));
defparam \fp_functions_0|expSum_uid44_fpMulTest_o[6] .is_wysiwyg = "true";
defparam \fp_functions_0|expSum_uid44_fpMulTest_o[6] .power_up = "low";

dffeas \fp_functions_0|expSum_uid44_fpMulTest_o[7] (
	.clk(clk),
	.d(\fp_functions_0|add_4~29_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|expSum_uid44_fpMulTest_o[7]~q ),
	.prn(vcc));
defparam \fp_functions_0|expSum_uid44_fpMulTest_o[7] .is_wysiwyg = "true";
defparam \fp_functions_0|expSum_uid44_fpMulTest_o[7] .power_up = "low";

dffeas \fp_functions_0|expSum_uid44_fpMulTest_o[8] (
	.clk(clk),
	.d(\fp_functions_0|add_4~33_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|expSum_uid44_fpMulTest_o[8]~q ),
	.prn(vcc));
defparam \fp_functions_0|expSum_uid44_fpMulTest_o[8] .is_wysiwyg = "true";
defparam \fp_functions_0|expSum_uid44_fpMulTest_o[8] .power_up = "low";

dffeas \fp_functions_0|expSum_uid44_fpMulTest_o[9] (
	.clk(clk),
	.d(\fp_functions_0|add_4~37_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|expSum_uid44_fpMulTest_o[9]~q ),
	.prn(vcc));
defparam \fp_functions_0|expSum_uid44_fpMulTest_o[9] .is_wysiwyg = "true";
defparam \fp_functions_0|expSum_uid44_fpMulTest_o[9] .power_up = "low";

dffeas \fp_functions_0|expSum_uid44_fpMulTest_o[10] (
	.clk(clk),
	.d(\fp_functions_0|add_4~41_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|expSum_uid44_fpMulTest_o[10]~q ),
	.prn(vcc));
defparam \fp_functions_0|expSum_uid44_fpMulTest_o[10] .is_wysiwyg = "true";
defparam \fp_functions_0|expSum_uid44_fpMulTest_o[10] .power_up = "low";

dffeas \fp_functions_0|signR_uid48_fpMulTest_delay|delay_signals[0][0] (
	.clk(clk),
	.d(\fp_functions_0|i1068~combout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|signR_uid48_fpMulTest_delay|delay_signals[0][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|signR_uid48_fpMulTest_delay|delay_signals[0][0] .is_wysiwyg = "true";
defparam \fp_functions_0|signR_uid48_fpMulTest_delay|delay_signals[0][0] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][0] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][0] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][0] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][1] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][1]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][1]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][1] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][1] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][2] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][2]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][2]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][2] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][2] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][3] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][3]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][3]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][3] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][3] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][4] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][4]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][4]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][4] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][4] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][5] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][5]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][5]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][5] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][5] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][6] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][6]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][6]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][6] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][6] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][7] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][7]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][7]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][7] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][7] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][8] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][8]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][8]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][8] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][8] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][9] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][9]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][9]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][9] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][9] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][10] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][10]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][10]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][10] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][10] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][11] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][11]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][11]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][11] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][11] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][12] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][12]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][12]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][12] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][12] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][13] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][13]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][13]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][13] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][13] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][14] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][14]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][14]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][14] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][14] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][15] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][15]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][15]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][15] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][15] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][16] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][16]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][16]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][16] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][16] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][17] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][17]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][17]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][17] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][17] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][18] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][18]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][18]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][18] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][18] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][19] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][19]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][19]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][19] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][19] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][20] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][20]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][20]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][20] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][20] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][21] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][21]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][21]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][21] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][21] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][22] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][22]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][22]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][22] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][22] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][23] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][23]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][23]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][23] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][23] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][24] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][24]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][24]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][24] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][24] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][25] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][25]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][25]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][25] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][25] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][26] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][26]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][26]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][26] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[0][26] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][0] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][0] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][0] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][1] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][1]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][1]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][1] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][1] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][2] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][2]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][2]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][2] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][2] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][3] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][3]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][3]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][3] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][3] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][4] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][4]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][4]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][4] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][4] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][5] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][5]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][5]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][5] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][5] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][6] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][6]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][6]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][6] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][6] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][7] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][7]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][7]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][7] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][7] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][8] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][8]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][8]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][8] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][8] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][9] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][9]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][9]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][9] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][9] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][10] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][10]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][10]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][10] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][10] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][11] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][11]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][11]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][11] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][11] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][12] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][12]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][12]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][12] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][12] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][13] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][13]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][13]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][13] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][13] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][14] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][14]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][14]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][14] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][14] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][15] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][15]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][15]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][15] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][15] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][16] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][16]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][16]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][16] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][16] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][17] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][17]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][17]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][17] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][17] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][18] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][18]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][18]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][18] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][18] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][19] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][19]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][19]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][19] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][19] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][20] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][20]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][20]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][20] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][20] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][21] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][21]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][21]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][21] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][21] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][22] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][22]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][22]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][22] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][22] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][23] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][23]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][23]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][23] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][23] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][24] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][24]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][24]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][24] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][24] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][25] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][25]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][25]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][25] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][25] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][26] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][26]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][26]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][26] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[0][26] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][0] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][0] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][0] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][1] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][1]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][1]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][1] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][1] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][2] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][2]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][2]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][2] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][2] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][3] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][3]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][3]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][3] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][3] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][4] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][4]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][4]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][4] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][4] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][5] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][5]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][5]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][5] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][5] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][6] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][6]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][6]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][6] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][6] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][7] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][7]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][7]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][7] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][7] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][8] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][8]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][8]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][8] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][8] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][9] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][9]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][9]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][9] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][9] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][10] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][10]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][10]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][10] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][10] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][11] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][11]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][11]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][11] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][11] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][12] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][12]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][12]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][12] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][12] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][13] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][13]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][13]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][13] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][13] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][14] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][14]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][14]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][14] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][14] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][15] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][15]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][15]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][15] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][15] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][16] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][16]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][16]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][16] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][16] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][17] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][17]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][17]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][17] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][17] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][18] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][18]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][18]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][18] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][18] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][19] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][19]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][19]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][19] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][19] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][20] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][20]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][20]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][20] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][20] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][21] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][21]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][21]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][21] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][21] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][22] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][22]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][22]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][22] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][22] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][23] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][23]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][23]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][23] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][23] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][24] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][24]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][24]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][24] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][24] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][25] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][25]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][25]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][25] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][25] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][26] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][26]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][26]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][26] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a1[0][26] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][0] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][0] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][0] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][1] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][1]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][1]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][1] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][1] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][2] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][2]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][2]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][2] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][2] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][3] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][3]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][3]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][3] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][3] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][4] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][4]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][4]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][4] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][4] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][5] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][5]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][5]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][5] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][5] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][6] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][6]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][6]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][6] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][6] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][7] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][7]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][7]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][7] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][7] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][8] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][8]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][8]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][8] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][8] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][9] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][9]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][9]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][9] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][9] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][10] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][10]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][10]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][10] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][10] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][11] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][11]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][11]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][11] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][11] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][12] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][12]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][12]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][12] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][12] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][13] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][13]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][13]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][13] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][13] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][14] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][14]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][14]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][14] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][14] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][15] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][15]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][15]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][15] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][15] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][16] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][16]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][16]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][16] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][16] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][17] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][17]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][17]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][17] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][17] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][18] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][18]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][18]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][18] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][18] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][19] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][19]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][19]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][19] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][19] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][20] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][20]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][20]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][20] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][20] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][21] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][21]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][21]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][21] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][21] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][22] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][22]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][22]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][22] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][22] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][23] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][23]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][23]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][23] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][23] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][24] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][24]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][24]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][24] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][24] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][25] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][25]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][25]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][25] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][25] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][26] (
	.clk(clk),
	.d(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][26]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][26]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][26] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c1[0][26] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][0] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][0] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][0] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][1] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][1]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][1]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][1] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][1] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][2] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][2]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][2]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][2] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][2] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][3] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][3]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][3]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][3] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][3] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][4] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][4]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][4]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][4] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][4] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][5] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][5]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][5]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][5] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][5] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][6] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][6]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][6]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][6] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][6] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][7] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][7]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][7]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][7] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][7] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][8] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][8]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][8]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][8] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][8] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][9] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][9]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][9]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][9] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][9] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][10] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][10]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][10]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][10] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][10] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][11] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][11]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][11]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][11] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][11] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][12] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][12]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][12]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][12] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][12] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][13] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][13]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][13]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][13] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][13] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][14] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][14]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][14]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][14] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][14] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][15] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][15]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][15]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][15] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][15] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][16] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][16]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][16]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][16] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][16] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][17] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][17]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][17]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][17] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][17] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][18] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][18]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][18]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][18] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][18] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][19] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][19]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][19]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][19] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][19] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][20] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][20]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][20]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][20] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][20] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][21] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][21]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][21]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][21] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][21] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][22] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][22]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][22]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][22] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][22] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][23] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][23]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][23]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][23] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][23] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][24] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][24]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][24]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][24] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][24] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][25] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][25]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][25]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][25] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][25] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][26] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][26]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][26]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][26] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a1[0][26] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][0] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][0] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][0] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][1] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][1]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][1]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][1] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][1] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][2] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][2]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][2]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][2] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][2] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][3] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][3]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][3]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][3] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][3] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][4] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][4]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][4]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][4] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][4] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][5] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][5]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][5]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][5] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][5] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][6] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][6]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][6]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][6] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][6] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][7] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][7]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][7]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][7] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][7] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][8] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][8]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][8]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][8] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][8] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][9] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][9]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][9]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][9] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][9] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][10] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][10]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][10]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][10] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][10] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][11] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][11]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][11]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][11] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][11] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][12] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][12]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][12]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][12] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][12] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][13] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][13]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][13]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][13] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][13] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][14] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][14]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][14]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][14] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][14] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][15] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][15]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][15]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][15] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][15] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][16] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][16]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][16]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][16] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][16] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][17] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][17]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][17]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][17] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][17] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][18] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][18]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][18]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][18] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][18] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][19] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][19]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][19]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][19] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][19] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][20] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][20]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][20]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][20] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][20] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][21] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][21]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][21]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][21] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][21] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][22] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][22]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][22]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][22] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][22] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][23] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][23]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][23]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][23] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][23] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][24] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][24]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][24]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][24] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][24] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][25] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][25]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][25]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][25] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][25] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][26] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][26]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][26]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][26] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c1[0][26] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|reduce_nor_2~0 (
	.dataa(!b[52]),
	.datab(!b[53]),
	.datac(!b[54]),
	.datad(!b[55]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|reduce_nor_2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|reduce_nor_2~0 .extended_lut = "off";
defparam \fp_functions_0|reduce_nor_2~0 .lut_mask = 64'h8000800080008000;
defparam \fp_functions_0|reduce_nor_2~0 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|reduce_nor_2~1 (
	.dataa(!b[58]),
	.datab(!b[59]),
	.datac(!b[60]),
	.datad(!b[61]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|reduce_nor_2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|reduce_nor_2~1 .extended_lut = "off";
defparam \fp_functions_0|reduce_nor_2~1 .lut_mask = 64'h8000800080008000;
defparam \fp_functions_0|reduce_nor_2~1 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|reduce_nor_2 (
	.dataa(!b[56]),
	.datab(!b[57]),
	.datac(!b[62]),
	.datad(!\fp_functions_0|reduce_nor_2~0_combout ),
	.datae(!\fp_functions_0|reduce_nor_2~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|reduce_nor_2~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|reduce_nor_2 .extended_lut = "off";
defparam \fp_functions_0|reduce_nor_2 .lut_mask = 64'h0000008000000080;
defparam \fp_functions_0|reduce_nor_2 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|reduce_nor_4~0 (
	.dataa(!b[52]),
	.datab(!b[53]),
	.datac(!b[54]),
	.datad(!b[55]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|reduce_nor_4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|reduce_nor_4~0 .extended_lut = "off";
defparam \fp_functions_0|reduce_nor_4~0 .lut_mask = 64'h0001000100010001;
defparam \fp_functions_0|reduce_nor_4~0 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|reduce_nor_4~1 (
	.dataa(!b[58]),
	.datab(!b[59]),
	.datac(!b[60]),
	.datad(!b[61]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|reduce_nor_4~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|reduce_nor_4~1 .extended_lut = "off";
defparam \fp_functions_0|reduce_nor_4~1 .lut_mask = 64'h0001000100010001;
defparam \fp_functions_0|reduce_nor_4~1 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|reduce_nor_4 (
	.dataa(!b[56]),
	.datab(!b[57]),
	.datac(!b[62]),
	.datad(!\fp_functions_0|reduce_nor_4~0_combout ),
	.datae(!\fp_functions_0|reduce_nor_4~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|reduce_nor_4~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|reduce_nor_4 .extended_lut = "off";
defparam \fp_functions_0|reduce_nor_4 .lut_mask = 64'h0000000100000001;
defparam \fp_functions_0|reduce_nor_4 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|reduce_nor_1~0 (
	.dataa(!a[52]),
	.datab(!a[53]),
	.datac(!a[54]),
	.datad(!a[55]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|reduce_nor_1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|reduce_nor_1~0 .extended_lut = "off";
defparam \fp_functions_0|reduce_nor_1~0 .lut_mask = 64'h0001000100010001;
defparam \fp_functions_0|reduce_nor_1~0 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|reduce_nor_1~1 (
	.dataa(!a[58]),
	.datab(!a[59]),
	.datac(!a[60]),
	.datad(!a[61]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|reduce_nor_1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|reduce_nor_1~1 .extended_lut = "off";
defparam \fp_functions_0|reduce_nor_1~1 .lut_mask = 64'h0001000100010001;
defparam \fp_functions_0|reduce_nor_1~1 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|reduce_nor_1 (
	.dataa(!a[56]),
	.datab(!a[57]),
	.datac(!a[62]),
	.datad(!\fp_functions_0|reduce_nor_1~0_combout ),
	.datae(!\fp_functions_0|reduce_nor_1~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|reduce_nor_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|reduce_nor_1 .extended_lut = "off";
defparam \fp_functions_0|reduce_nor_1 .lut_mask = 64'h0000000100000001;
defparam \fp_functions_0|reduce_nor_1 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|reduce_nor_5~0 (
	.dataa(!a[52]),
	.datab(!a[53]),
	.datac(!a[54]),
	.datad(!a[55]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|reduce_nor_5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|reduce_nor_5~0 .extended_lut = "off";
defparam \fp_functions_0|reduce_nor_5~0 .lut_mask = 64'h8000800080008000;
defparam \fp_functions_0|reduce_nor_5~0 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|reduce_nor_5~1 (
	.dataa(!a[58]),
	.datab(!a[59]),
	.datac(!a[60]),
	.datad(!a[61]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|reduce_nor_5~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|reduce_nor_5~1 .extended_lut = "off";
defparam \fp_functions_0|reduce_nor_5~1 .lut_mask = 64'h8000800080008000;
defparam \fp_functions_0|reduce_nor_5~1 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|reduce_nor_5 (
	.dataa(!a[56]),
	.datab(!a[57]),
	.datac(!a[62]),
	.datad(!\fp_functions_0|reduce_nor_5~0_combout ),
	.datae(!\fp_functions_0|reduce_nor_5~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|reduce_nor_5~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|reduce_nor_5 .extended_lut = "off";
defparam \fp_functions_0|reduce_nor_5 .lut_mask = 64'h0000008000000080;
defparam \fp_functions_0|reduce_nor_5 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|reduce_nor_3~0 (
	.dataa(!b[18]),
	.datab(!b[19]),
	.datac(!b[20]),
	.datad(!b[21]),
	.datae(!b[22]),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|reduce_nor_3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|reduce_nor_3~0 .extended_lut = "off";
defparam \fp_functions_0|reduce_nor_3~0 .lut_mask = 64'h8000000080000000;
defparam \fp_functions_0|reduce_nor_3~0 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|reduce_nor_3~1 (
	.dataa(!b[24]),
	.datab(!b[25]),
	.datac(!b[26]),
	.datad(!b[27]),
	.datae(!b[28]),
	.dataf(!b[29]),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|reduce_nor_3~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|reduce_nor_3~1 .extended_lut = "off";
defparam \fp_functions_0|reduce_nor_3~1 .lut_mask = 64'h8000000000000000;
defparam \fp_functions_0|reduce_nor_3~1 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|reduce_nor_3~2 (
	.dataa(!b[30]),
	.datab(!b[31]),
	.datac(!b[32]),
	.datad(!b[33]),
	.datae(!b[34]),
	.dataf(!b[35]),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|reduce_nor_3~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|reduce_nor_3~2 .extended_lut = "off";
defparam \fp_functions_0|reduce_nor_3~2 .lut_mask = 64'h8000000000000000;
defparam \fp_functions_0|reduce_nor_3~2 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|reduce_nor_3~3 (
	.dataa(!b[0]),
	.datab(!b[1]),
	.datac(!b[2]),
	.datad(!b[3]),
	.datae(!b[4]),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|reduce_nor_3~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|reduce_nor_3~3 .extended_lut = "off";
defparam \fp_functions_0|reduce_nor_3~3 .lut_mask = 64'h8000000080000000;
defparam \fp_functions_0|reduce_nor_3~3 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|reduce_nor_3~4 (
	.dataa(!b[6]),
	.datab(!b[7]),
	.datac(!b[8]),
	.datad(!b[9]),
	.datae(!b[10]),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|reduce_nor_3~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|reduce_nor_3~4 .extended_lut = "off";
defparam \fp_functions_0|reduce_nor_3~4 .lut_mask = 64'h8000000080000000;
defparam \fp_functions_0|reduce_nor_3~4 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|reduce_nor_3~5 (
	.dataa(!b[12]),
	.datab(!b[13]),
	.datac(!b[14]),
	.datad(!b[15]),
	.datae(!b[16]),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|reduce_nor_3~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|reduce_nor_3~5 .extended_lut = "off";
defparam \fp_functions_0|reduce_nor_3~5 .lut_mask = 64'h8000000080000000;
defparam \fp_functions_0|reduce_nor_3~5 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|reduce_nor_3~6 (
	.dataa(!b[5]),
	.datab(!b[11]),
	.datac(!b[17]),
	.datad(!\fp_functions_0|reduce_nor_3~3_combout ),
	.datae(!\fp_functions_0|reduce_nor_3~4_combout ),
	.dataf(!\fp_functions_0|reduce_nor_3~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|reduce_nor_3~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|reduce_nor_3~6 .extended_lut = "off";
defparam \fp_functions_0|reduce_nor_3~6 .lut_mask = 64'h0000000000000080;
defparam \fp_functions_0|reduce_nor_3~6 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|reduce_nor_3~7 (
	.dataa(!b[48]),
	.datab(!b[49]),
	.datac(!b[50]),
	.datad(!b[51]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|reduce_nor_3~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|reduce_nor_3~7 .extended_lut = "off";
defparam \fp_functions_0|reduce_nor_3~7 .lut_mask = 64'h8000800080008000;
defparam \fp_functions_0|reduce_nor_3~7 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|reduce_nor_3~8 (
	.dataa(!b[36]),
	.datab(!b[37]),
	.datac(!b[38]),
	.datad(!b[39]),
	.datae(!b[40]),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|reduce_nor_3~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|reduce_nor_3~8 .extended_lut = "off";
defparam \fp_functions_0|reduce_nor_3~8 .lut_mask = 64'h8000000080000000;
defparam \fp_functions_0|reduce_nor_3~8 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|reduce_nor_3~9 (
	.dataa(!b[42]),
	.datab(!b[43]),
	.datac(!b[44]),
	.datad(!b[45]),
	.datae(!b[46]),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|reduce_nor_3~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|reduce_nor_3~9 .extended_lut = "off";
defparam \fp_functions_0|reduce_nor_3~9 .lut_mask = 64'h8000000080000000;
defparam \fp_functions_0|reduce_nor_3~9 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|reduce_nor_3~10 (
	.dataa(!b[41]),
	.datab(!b[47]),
	.datac(!\fp_functions_0|reduce_nor_3~7_combout ),
	.datad(!\fp_functions_0|reduce_nor_3~8_combout ),
	.datae(!\fp_functions_0|reduce_nor_3~9_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|reduce_nor_3~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|reduce_nor_3~10 .extended_lut = "off";
defparam \fp_functions_0|reduce_nor_3~10 .lut_mask = 64'h0000000800000008;
defparam \fp_functions_0|reduce_nor_3~10 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|reduce_nor_3 (
	.dataa(!b[23]),
	.datab(!\fp_functions_0|reduce_nor_3~0_combout ),
	.datac(!\fp_functions_0|reduce_nor_3~1_combout ),
	.datad(!\fp_functions_0|reduce_nor_3~2_combout ),
	.datae(!\fp_functions_0|reduce_nor_3~6_combout ),
	.dataf(!\fp_functions_0|reduce_nor_3~10_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|reduce_nor_3~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|reduce_nor_3 .extended_lut = "off";
defparam \fp_functions_0|reduce_nor_3 .lut_mask = 64'h0000000000000002;
defparam \fp_functions_0|reduce_nor_3 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|reduce_nor_0~0 (
	.dataa(!a[18]),
	.datab(!a[19]),
	.datac(!a[20]),
	.datad(!a[21]),
	.datae(!a[22]),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|reduce_nor_0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|reduce_nor_0~0 .extended_lut = "off";
defparam \fp_functions_0|reduce_nor_0~0 .lut_mask = 64'h8000000080000000;
defparam \fp_functions_0|reduce_nor_0~0 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|reduce_nor_0~1 (
	.dataa(!a[24]),
	.datab(!a[25]),
	.datac(!a[26]),
	.datad(!a[27]),
	.datae(!a[28]),
	.dataf(!a[29]),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|reduce_nor_0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|reduce_nor_0~1 .extended_lut = "off";
defparam \fp_functions_0|reduce_nor_0~1 .lut_mask = 64'h8000000000000000;
defparam \fp_functions_0|reduce_nor_0~1 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|reduce_nor_0~2 (
	.dataa(!a[30]),
	.datab(!a[31]),
	.datac(!a[32]),
	.datad(!a[33]),
	.datae(!a[34]),
	.dataf(!a[35]),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|reduce_nor_0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|reduce_nor_0~2 .extended_lut = "off";
defparam \fp_functions_0|reduce_nor_0~2 .lut_mask = 64'h8000000000000000;
defparam \fp_functions_0|reduce_nor_0~2 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|reduce_nor_0~3 (
	.dataa(!a[0]),
	.datab(!a[1]),
	.datac(!a[2]),
	.datad(!a[3]),
	.datae(!a[4]),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|reduce_nor_0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|reduce_nor_0~3 .extended_lut = "off";
defparam \fp_functions_0|reduce_nor_0~3 .lut_mask = 64'h8000000080000000;
defparam \fp_functions_0|reduce_nor_0~3 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|reduce_nor_0~4 (
	.dataa(!a[6]),
	.datab(!a[7]),
	.datac(!a[8]),
	.datad(!a[9]),
	.datae(!a[10]),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|reduce_nor_0~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|reduce_nor_0~4 .extended_lut = "off";
defparam \fp_functions_0|reduce_nor_0~4 .lut_mask = 64'h8000000080000000;
defparam \fp_functions_0|reduce_nor_0~4 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|reduce_nor_0~5 (
	.dataa(!a[12]),
	.datab(!a[13]),
	.datac(!a[14]),
	.datad(!a[15]),
	.datae(!a[16]),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|reduce_nor_0~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|reduce_nor_0~5 .extended_lut = "off";
defparam \fp_functions_0|reduce_nor_0~5 .lut_mask = 64'h8000000080000000;
defparam \fp_functions_0|reduce_nor_0~5 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|reduce_nor_0~6 (
	.dataa(!a[5]),
	.datab(!a[11]),
	.datac(!a[17]),
	.datad(!\fp_functions_0|reduce_nor_0~3_combout ),
	.datae(!\fp_functions_0|reduce_nor_0~4_combout ),
	.dataf(!\fp_functions_0|reduce_nor_0~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|reduce_nor_0~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|reduce_nor_0~6 .extended_lut = "off";
defparam \fp_functions_0|reduce_nor_0~6 .lut_mask = 64'h0000000000000080;
defparam \fp_functions_0|reduce_nor_0~6 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|reduce_nor_0~7 (
	.dataa(!a[48]),
	.datab(!a[49]),
	.datac(!a[50]),
	.datad(!a[51]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|reduce_nor_0~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|reduce_nor_0~7 .extended_lut = "off";
defparam \fp_functions_0|reduce_nor_0~7 .lut_mask = 64'h8000800080008000;
defparam \fp_functions_0|reduce_nor_0~7 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|reduce_nor_0~8 (
	.dataa(!a[36]),
	.datab(!a[37]),
	.datac(!a[38]),
	.datad(!a[39]),
	.datae(!a[40]),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|reduce_nor_0~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|reduce_nor_0~8 .extended_lut = "off";
defparam \fp_functions_0|reduce_nor_0~8 .lut_mask = 64'h8000000080000000;
defparam \fp_functions_0|reduce_nor_0~8 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|reduce_nor_0~9 (
	.dataa(!a[42]),
	.datab(!a[43]),
	.datac(!a[44]),
	.datad(!a[45]),
	.datae(!a[46]),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|reduce_nor_0~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|reduce_nor_0~9 .extended_lut = "off";
defparam \fp_functions_0|reduce_nor_0~9 .lut_mask = 64'h8000000080000000;
defparam \fp_functions_0|reduce_nor_0~9 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|reduce_nor_0~10 (
	.dataa(!a[41]),
	.datab(!a[47]),
	.datac(!\fp_functions_0|reduce_nor_0~7_combout ),
	.datad(!\fp_functions_0|reduce_nor_0~8_combout ),
	.datae(!\fp_functions_0|reduce_nor_0~9_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|reduce_nor_0~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|reduce_nor_0~10 .extended_lut = "off";
defparam \fp_functions_0|reduce_nor_0~10 .lut_mask = 64'h0000000800000008;
defparam \fp_functions_0|reduce_nor_0~10 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|reduce_nor_0 (
	.dataa(!a[23]),
	.datab(!\fp_functions_0|reduce_nor_0~0_combout ),
	.datac(!\fp_functions_0|reduce_nor_0~1_combout ),
	.datad(!\fp_functions_0|reduce_nor_0~2_combout ),
	.datae(!\fp_functions_0|reduce_nor_0~6_combout ),
	.dataf(!\fp_functions_0|reduce_nor_0~10_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|reduce_nor_0~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|reduce_nor_0 .extended_lut = "off";
defparam \fp_functions_0|reduce_nor_0 .lut_mask = 64'h0000000000000002;
defparam \fp_functions_0|reduce_nor_0 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|reduce_nor_9 (
	.dataa(!\fp_functions_0|redist15_rdcnt_i[0]~q ),
	.datab(!\fp_functions_0|redist15_rdcnt_i[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|reduce_nor_9~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|reduce_nor_9 .extended_lut = "off";
defparam \fp_functions_0|reduce_nor_9 .lut_mask = 64'h8888888888888888;
defparam \fp_functions_0|reduce_nor_9 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|i1068 (
	.dataa(!a[63]),
	.datab(!b[63]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|i1068~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|i1068 .extended_lut = "off";
defparam \fp_functions_0|i1068 .lut_mask = 64'h6666666666666666;
defparam \fp_functions_0|i1068 .shared_arith = "off";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][0] (
	.clk(clk),
	.d(\fp_functions_0|redist6|delay_signals[0][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][0] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][0] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][1] (
	.clk(clk),
	.d(\fp_functions_0|redist6|delay_signals[0][1]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][1]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][1] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][1] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][2] (
	.clk(clk),
	.d(\fp_functions_0|redist6|delay_signals[0][2]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][2]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][2] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][2] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][3] (
	.clk(clk),
	.d(\fp_functions_0|redist6|delay_signals[0][3]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][3]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][3] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][3] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][4] (
	.clk(clk),
	.d(\fp_functions_0|redist6|delay_signals[0][4]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][4]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][4] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][4] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][5] (
	.clk(clk),
	.d(\fp_functions_0|redist6|delay_signals[0][5]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][5]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][5] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][5] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][6] (
	.clk(clk),
	.d(\fp_functions_0|redist6|delay_signals[0][6]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][6]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][6] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][6] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][7] (
	.clk(clk),
	.d(\fp_functions_0|redist6|delay_signals[0][7]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][7]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][7] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][7] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][8] (
	.clk(clk),
	.d(\fp_functions_0|redist6|delay_signals[0][8]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][8]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][8] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][8] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][9] (
	.clk(clk),
	.d(\fp_functions_0|redist6|delay_signals[0][9]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][9]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][9] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][9] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][10] (
	.clk(clk),
	.d(\fp_functions_0|redist6|delay_signals[0][10]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][10]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][10] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][10] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][11] (
	.clk(clk),
	.d(\fp_functions_0|redist6|delay_signals[0][11]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][11]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][11] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][11] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][12] (
	.clk(clk),
	.d(\fp_functions_0|redist6|delay_signals[0][12]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][12]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][12] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][12] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][13] (
	.clk(clk),
	.d(\fp_functions_0|redist6|delay_signals[0][13]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][13]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][13] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][13] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][14] (
	.clk(clk),
	.d(\fp_functions_0|redist6|delay_signals[0][14]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][14]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][14] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][14] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][15] (
	.clk(clk),
	.d(\fp_functions_0|redist6|delay_signals[0][15]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][15]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][15] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][15] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][16] (
	.clk(clk),
	.d(\fp_functions_0|redist6|delay_signals[0][16]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][16]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][16] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][16] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][17] (
	.clk(clk),
	.d(\fp_functions_0|redist6|delay_signals[0][17]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][17]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][17] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][17] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][18] (
	.clk(clk),
	.d(\fp_functions_0|redist6|delay_signals[0][18]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][18]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][18] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][18] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][19] (
	.clk(clk),
	.d(\fp_functions_0|redist6|delay_signals[0][19]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][19]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][19] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][19] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][20] (
	.clk(clk),
	.d(\fp_functions_0|redist6|delay_signals[0][20]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][20]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][20] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][20] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][21] (
	.clk(clk),
	.d(\fp_functions_0|redist6|delay_signals[0][21]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][21]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][21] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][21] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][22] (
	.clk(clk),
	.d(\fp_functions_0|redist6|delay_signals[0][22]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][22]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][22] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][22] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][23] (
	.clk(clk),
	.d(\fp_functions_0|redist6|delay_signals[0][23]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][23]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][23] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][23] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][24] (
	.clk(clk),
	.d(\fp_functions_0|redist6|delay_signals[0][24]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][24]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][24] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][24] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][25] (
	.clk(clk),
	.d(\fp_functions_0|redist6|delay_signals[0][25]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][25]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][25] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][25] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][26] (
	.clk(clk),
	.d(\fp_functions_0|redist6|delay_signals[0][26]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][26]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][26] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[0][26] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][0] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][0]~0_combout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][0] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][0] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][1] (
	.clk(clk),
	.d(\fp_functions_0|redist4|delay_signals[0][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][1]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][1] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][1] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][2] (
	.clk(clk),
	.d(\fp_functions_0|redist4|delay_signals[0][1]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][2]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][2] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][2] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][3] (
	.clk(clk),
	.d(\fp_functions_0|redist4|delay_signals[0][2]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][3]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][3] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][3] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][4] (
	.clk(clk),
	.d(\fp_functions_0|redist4|delay_signals[0][3]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][4]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][4] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][4] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][5] (
	.clk(clk),
	.d(\fp_functions_0|redist4|delay_signals[0][4]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][5]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][5] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][5] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][6] (
	.clk(clk),
	.d(\fp_functions_0|redist4|delay_signals[0][5]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][6]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][6] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][6] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][7] (
	.clk(clk),
	.d(\fp_functions_0|redist4|delay_signals[0][6]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][7]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][7] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][7] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][8] (
	.clk(clk),
	.d(\fp_functions_0|redist4|delay_signals[0][7]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][8]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][8] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][8] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][9] (
	.clk(clk),
	.d(\fp_functions_0|redist4|delay_signals[0][8]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][9]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][9] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][9] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][10] (
	.clk(clk),
	.d(\fp_functions_0|redist4|delay_signals[0][9]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][10]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][10] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][10] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][11] (
	.clk(clk),
	.d(\fp_functions_0|redist4|delay_signals[0][10]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][11]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][11] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][11] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][12] (
	.clk(clk),
	.d(\fp_functions_0|redist4|delay_signals[0][11]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][12]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][12] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][12] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][13] (
	.clk(clk),
	.d(\fp_functions_0|redist4|delay_signals[0][12]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][13]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][13] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][13] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][14] (
	.clk(clk),
	.d(\fp_functions_0|redist4|delay_signals[0][13]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][14]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][14] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][14] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][15] (
	.clk(clk),
	.d(\fp_functions_0|redist4|delay_signals[0][14]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][15]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][15] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][15] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][16] (
	.clk(clk),
	.d(\fp_functions_0|redist4|delay_signals[0][15]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][16]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][16] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][16] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][17] (
	.clk(clk),
	.d(\fp_functions_0|redist4|delay_signals[0][16]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][17]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][17] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][17] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][18] (
	.clk(clk),
	.d(\fp_functions_0|redist4|delay_signals[0][17]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][18]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][18] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][18] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][19] (
	.clk(clk),
	.d(\fp_functions_0|redist4|delay_signals[0][18]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][19]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][19] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][19] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][20] (
	.clk(clk),
	.d(\fp_functions_0|redist4|delay_signals[0][19]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][20]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][20] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][20] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][21] (
	.clk(clk),
	.d(\fp_functions_0|redist4|delay_signals[0][20]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][21]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][21] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][21] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][22] (
	.clk(clk),
	.d(\fp_functions_0|redist4|delay_signals[0][21]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][22]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][22] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][22] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][23] (
	.clk(clk),
	.d(\fp_functions_0|redist4|delay_signals[0][22]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][23]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][23] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][23] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][24] (
	.clk(clk),
	.d(\fp_functions_0|redist4|delay_signals[0][23]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][24]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][24] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][24] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][25] (
	.clk(clk),
	.d(\fp_functions_0|redist4|delay_signals[0][24]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][25]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][25] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][25] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][26] (
	.clk(clk),
	.d(\fp_functions_0|redist4|delay_signals[0][25]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][26]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][26] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][26] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][0] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][0] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][0] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][1] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][1]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][1]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][1] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][1] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][2] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][2]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][2]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][2] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][2] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][3] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][3]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][3]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][3] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][3] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][4] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][4]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][4]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][4] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][4] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][5] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][5]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][5]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][5] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][5] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][6] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][6]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][6]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][6] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][6] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][7] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][7]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][7]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][7] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][7] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][8] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][8]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][8]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][8] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][8] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][9] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][9]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][9]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][9] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][9] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][10] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][10]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][10]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][10] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][10] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][11] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][11]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][11]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][11] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][11] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][12] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][12]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][12]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][12] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][12] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][13] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][13]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][13]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][13] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][13] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][14] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][14]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][14]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][14] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][14] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][15] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][15]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][15]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][15] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][15] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][16] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][16]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][16]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][16] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][16] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][17] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][17]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][17]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][17] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][17] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][18] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][18]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][18]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][18] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][18] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][19] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][19]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][19]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][19] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][19] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][20] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][20]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][20]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][20] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][20] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][21] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][21]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][21]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][21] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][21] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][22] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][22]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][22]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][22] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][22] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][23] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][23]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][23]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][23] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][23] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][24] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][24]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][24]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][24] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][24] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][25] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][25]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][25]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][25] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][25] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][26] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][26]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][26]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][26] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a1[1][26] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][0] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][0] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][0] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][1] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][1]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][1]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][1] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][1] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][2] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][2]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][2]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][2] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][2] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][3] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][3]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][3]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][3] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][3] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][4] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][4]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][4]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][4] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][4] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][5] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][5]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][5]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][5] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][5] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][6] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][6]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][6]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][6] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][6] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][7] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][7]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][7]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][7] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][7] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][8] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][8]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][8]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][8] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][8] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][9] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][9]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][9]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][9] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][9] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][10] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][10]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][10]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][10] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][10] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][11] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][11]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][11]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][11] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][11] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][12] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][12]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][12]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][12] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][12] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][13] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][13]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][13]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][13] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][13] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][14] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][14]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][14]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][14] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][14] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][15] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][15]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][15]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][15] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][15] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][16] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][16]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][16]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][16] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][16] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][17] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][17]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][17]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][17] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][17] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][18] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][18]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][18]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][18] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][18] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][19] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][19]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][19]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][19] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][19] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][20] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][20]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][20]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][20] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][20] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][21] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][21]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][21]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][21] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][21] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][22] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][22]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][22]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][22] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][22] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][23] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][23]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][23]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][23] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][23] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][24] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][24]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][24]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][24] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][24] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][25] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][25]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][25]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][25] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][25] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][26] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][26]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][26]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][26] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c1[1][26] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][0] (
	.clk(clk),
	.d(\fp_functions_0|redist7|delay_signals[0][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][0] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][0] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][1] (
	.clk(clk),
	.d(\fp_functions_0|redist7|delay_signals[0][1]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][1]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][1] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][1] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][2] (
	.clk(clk),
	.d(\fp_functions_0|redist7|delay_signals[0][2]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][2]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][2] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][2] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][3] (
	.clk(clk),
	.d(\fp_functions_0|redist7|delay_signals[0][3]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][3]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][3] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][3] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][4] (
	.clk(clk),
	.d(\fp_functions_0|redist7|delay_signals[0][4]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][4]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][4] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][4] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][5] (
	.clk(clk),
	.d(\fp_functions_0|redist7|delay_signals[0][5]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][5]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][5] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][5] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][6] (
	.clk(clk),
	.d(\fp_functions_0|redist7|delay_signals[0][6]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][6]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][6] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][6] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][7] (
	.clk(clk),
	.d(\fp_functions_0|redist7|delay_signals[0][7]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][7]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][7] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][7] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][8] (
	.clk(clk),
	.d(\fp_functions_0|redist7|delay_signals[0][8]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][8]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][8] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][8] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][9] (
	.clk(clk),
	.d(\fp_functions_0|redist7|delay_signals[0][9]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][9]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][9] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][9] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][10] (
	.clk(clk),
	.d(\fp_functions_0|redist7|delay_signals[0][10]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][10]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][10] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][10] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][11] (
	.clk(clk),
	.d(\fp_functions_0|redist7|delay_signals[0][11]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][11]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][11] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][11] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][12] (
	.clk(clk),
	.d(\fp_functions_0|redist7|delay_signals[0][12]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][12]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][12] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][12] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][13] (
	.clk(clk),
	.d(\fp_functions_0|redist7|delay_signals[0][13]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][13]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][13] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][13] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][14] (
	.clk(clk),
	.d(\fp_functions_0|redist7|delay_signals[0][14]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][14]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][14] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][14] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][15] (
	.clk(clk),
	.d(\fp_functions_0|redist7|delay_signals[0][15]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][15]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][15] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][15] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][16] (
	.clk(clk),
	.d(\fp_functions_0|redist7|delay_signals[0][16]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][16]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][16] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][16] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][17] (
	.clk(clk),
	.d(\fp_functions_0|redist7|delay_signals[0][17]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][17]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][17] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][17] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][18] (
	.clk(clk),
	.d(\fp_functions_0|redist7|delay_signals[0][18]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][18]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][18] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][18] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][19] (
	.clk(clk),
	.d(\fp_functions_0|redist7|delay_signals[0][19]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][19]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][19] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][19] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][20] (
	.clk(clk),
	.d(\fp_functions_0|redist7|delay_signals[0][20]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][20]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][20] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][20] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][21] (
	.clk(clk),
	.d(\fp_functions_0|redist7|delay_signals[0][21]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][21]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][21] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][21] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][22] (
	.clk(clk),
	.d(\fp_functions_0|redist7|delay_signals[0][22]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][22]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][22] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][22] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][23] (
	.clk(clk),
	.d(\fp_functions_0|redist7|delay_signals[0][23]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][23]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][23] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][23] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][24] (
	.clk(clk),
	.d(\fp_functions_0|redist7|delay_signals[0][24]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][24]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][24] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][24] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][25] (
	.clk(clk),
	.d(\fp_functions_0|redist7|delay_signals[0][25]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][25]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][25] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][25] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][26] (
	.clk(clk),
	.d(\fp_functions_0|redist7|delay_signals[0][26]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][26]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][26] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_a0[0][26] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][0] (
	.clk(clk),
	.d(\fp_functions_0|redist6|delay_signals[0][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][0] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][0] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][1] (
	.clk(clk),
	.d(\fp_functions_0|redist6|delay_signals[0][1]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][1]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][1] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][1] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][2] (
	.clk(clk),
	.d(\fp_functions_0|redist6|delay_signals[0][2]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][2]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][2] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][2] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][3] (
	.clk(clk),
	.d(\fp_functions_0|redist6|delay_signals[0][3]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][3]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][3] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][3] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][4] (
	.clk(clk),
	.d(\fp_functions_0|redist6|delay_signals[0][4]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][4]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][4] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][4] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][5] (
	.clk(clk),
	.d(\fp_functions_0|redist6|delay_signals[0][5]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][5]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][5] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][5] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][6] (
	.clk(clk),
	.d(\fp_functions_0|redist6|delay_signals[0][6]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][6]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][6] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][6] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][7] (
	.clk(clk),
	.d(\fp_functions_0|redist6|delay_signals[0][7]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][7]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][7] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][7] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][8] (
	.clk(clk),
	.d(\fp_functions_0|redist6|delay_signals[0][8]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][8]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][8] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][8] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][9] (
	.clk(clk),
	.d(\fp_functions_0|redist6|delay_signals[0][9]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][9]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][9] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][9] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][10] (
	.clk(clk),
	.d(\fp_functions_0|redist6|delay_signals[0][10]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][10]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][10] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][10] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][11] (
	.clk(clk),
	.d(\fp_functions_0|redist6|delay_signals[0][11]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][11]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][11] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][11] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][12] (
	.clk(clk),
	.d(\fp_functions_0|redist6|delay_signals[0][12]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][12]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][12] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][12] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][13] (
	.clk(clk),
	.d(\fp_functions_0|redist6|delay_signals[0][13]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][13]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][13] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][13] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][14] (
	.clk(clk),
	.d(\fp_functions_0|redist6|delay_signals[0][14]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][14]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][14] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][14] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][15] (
	.clk(clk),
	.d(\fp_functions_0|redist6|delay_signals[0][15]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][15]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][15] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][15] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][16] (
	.clk(clk),
	.d(\fp_functions_0|redist6|delay_signals[0][16]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][16]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][16] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][16] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][17] (
	.clk(clk),
	.d(\fp_functions_0|redist6|delay_signals[0][17]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][17]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][17] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][17] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][18] (
	.clk(clk),
	.d(\fp_functions_0|redist6|delay_signals[0][18]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][18]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][18] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][18] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][19] (
	.clk(clk),
	.d(\fp_functions_0|redist6|delay_signals[0][19]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][19]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][19] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][19] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][20] (
	.clk(clk),
	.d(\fp_functions_0|redist6|delay_signals[0][20]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][20]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][20] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][20] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][21] (
	.clk(clk),
	.d(\fp_functions_0|redist6|delay_signals[0][21]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][21]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][21] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][21] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][22] (
	.clk(clk),
	.d(\fp_functions_0|redist6|delay_signals[0][22]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][22]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][22] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][22] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][23] (
	.clk(clk),
	.d(\fp_functions_0|redist6|delay_signals[0][23]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][23]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][23] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][23] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][24] (
	.clk(clk),
	.d(\fp_functions_0|redist6|delay_signals[0][24]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][24]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][24] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][24] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][25] (
	.clk(clk),
	.d(\fp_functions_0|redist6|delay_signals[0][25]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][25]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][25] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][25] .power_up = "low";

dffeas \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][26] (
	.clk(clk),
	.d(\fp_functions_0|redist6|delay_signals[0][26]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][26]~q ),
	.prn(vcc));
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][26] .is_wysiwyg = "true";
defparam \fp_functions_0|topProd_uid107_prod_uid47_fpMulTest_cma_c0[0][26] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][0] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][0]~0_combout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][0] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][0] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][1] (
	.clk(clk),
	.d(\fp_functions_0|redist4|delay_signals[0][0]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][1]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][1] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][1] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][2] (
	.clk(clk),
	.d(\fp_functions_0|redist4|delay_signals[0][1]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][2]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][2] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][2] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][3] (
	.clk(clk),
	.d(\fp_functions_0|redist4|delay_signals[0][2]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][3]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][3] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][3] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][4] (
	.clk(clk),
	.d(\fp_functions_0|redist4|delay_signals[0][3]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][4]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][4] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][4] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][5] (
	.clk(clk),
	.d(\fp_functions_0|redist4|delay_signals[0][4]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][5]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][5] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][5] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][6] (
	.clk(clk),
	.d(\fp_functions_0|redist4|delay_signals[0][5]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][6]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][6] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][6] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][7] (
	.clk(clk),
	.d(\fp_functions_0|redist4|delay_signals[0][6]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][7]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][7] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][7] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][8] (
	.clk(clk),
	.d(\fp_functions_0|redist4|delay_signals[0][7]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][8]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][8] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][8] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][9] (
	.clk(clk),
	.d(\fp_functions_0|redist4|delay_signals[0][8]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][9]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][9] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][9] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][10] (
	.clk(clk),
	.d(\fp_functions_0|redist4|delay_signals[0][9]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][10]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][10] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][10] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][11] (
	.clk(clk),
	.d(\fp_functions_0|redist4|delay_signals[0][10]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][11]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][11] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][11] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][12] (
	.clk(clk),
	.d(\fp_functions_0|redist4|delay_signals[0][11]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][12]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][12] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][12] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][13] (
	.clk(clk),
	.d(\fp_functions_0|redist4|delay_signals[0][12]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][13]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][13] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][13] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][14] (
	.clk(clk),
	.d(\fp_functions_0|redist4|delay_signals[0][13]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][14]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][14] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][14] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][15] (
	.clk(clk),
	.d(\fp_functions_0|redist4|delay_signals[0][14]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][15]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][15] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][15] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][16] (
	.clk(clk),
	.d(\fp_functions_0|redist4|delay_signals[0][15]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][16]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][16] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][16] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][17] (
	.clk(clk),
	.d(\fp_functions_0|redist4|delay_signals[0][16]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][17]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][17] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][17] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][18] (
	.clk(clk),
	.d(\fp_functions_0|redist4|delay_signals[0][17]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][18]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][18] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][18] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][19] (
	.clk(clk),
	.d(\fp_functions_0|redist4|delay_signals[0][18]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][19]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][19] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][19] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][20] (
	.clk(clk),
	.d(\fp_functions_0|redist4|delay_signals[0][19]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][20]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][20] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][20] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][21] (
	.clk(clk),
	.d(\fp_functions_0|redist4|delay_signals[0][20]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][21]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][21] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][21] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][22] (
	.clk(clk),
	.d(\fp_functions_0|redist4|delay_signals[0][21]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][22]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][22] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][22] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][23] (
	.clk(clk),
	.d(\fp_functions_0|redist4|delay_signals[0][22]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][23]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][23] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][23] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][24] (
	.clk(clk),
	.d(\fp_functions_0|redist4|delay_signals[0][23]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][24]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][24] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][24] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][25] (
	.clk(clk),
	.d(\fp_functions_0|redist4|delay_signals[0][24]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][25]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][25] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][25] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][26] (
	.clk(clk),
	.d(\fp_functions_0|redist4|delay_signals[0][25]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][26]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][26] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][26] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][0] (
	.clk(clk),
	.d(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][0]~0_combout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][0] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][0] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][1] (
	.clk(clk),
	.d(\fp_functions_0|redist5|delay_signals[0][1]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][1]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][1] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][1] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][2] (
	.clk(clk),
	.d(\fp_functions_0|redist5|delay_signals[0][2]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][2]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][2] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][2] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][3] (
	.clk(clk),
	.d(\fp_functions_0|redist5|delay_signals[0][3]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][3]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][3] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][3] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][4] (
	.clk(clk),
	.d(\fp_functions_0|redist5|delay_signals[0][4]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][4]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][4] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][4] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][5] (
	.clk(clk),
	.d(\fp_functions_0|redist5|delay_signals[0][5]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][5]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][5] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][5] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][6] (
	.clk(clk),
	.d(\fp_functions_0|redist5|delay_signals[0][6]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][6]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][6] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][6] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][7] (
	.clk(clk),
	.d(\fp_functions_0|redist5|delay_signals[0][7]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][7]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][7] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][7] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][8] (
	.clk(clk),
	.d(\fp_functions_0|redist5|delay_signals[0][8]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][8]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][8] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][8] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][9] (
	.clk(clk),
	.d(\fp_functions_0|redist5|delay_signals[0][9]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][9]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][9] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][9] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][10] (
	.clk(clk),
	.d(\fp_functions_0|redist5|delay_signals[0][10]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][10]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][10] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][10] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][11] (
	.clk(clk),
	.d(\fp_functions_0|redist5|delay_signals[0][11]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][11]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][11] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][11] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][12] (
	.clk(clk),
	.d(\fp_functions_0|redist5|delay_signals[0][12]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][12]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][12] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][12] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][13] (
	.clk(clk),
	.d(\fp_functions_0|redist5|delay_signals[0][13]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][13]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][13] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][13] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][14] (
	.clk(clk),
	.d(\fp_functions_0|redist5|delay_signals[0][14]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][14]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][14] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][14] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][15] (
	.clk(clk),
	.d(\fp_functions_0|redist5|delay_signals[0][15]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][15]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][15] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][15] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][16] (
	.clk(clk),
	.d(\fp_functions_0|redist5|delay_signals[0][16]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][16]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][16] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][16] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][17] (
	.clk(clk),
	.d(\fp_functions_0|redist5|delay_signals[0][17]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][17]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][17] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][17] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][18] (
	.clk(clk),
	.d(\fp_functions_0|redist5|delay_signals[0][18]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][18]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][18] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][18] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][19] (
	.clk(clk),
	.d(\fp_functions_0|redist5|delay_signals[0][19]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][19]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][19] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][19] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][20] (
	.clk(clk),
	.d(\fp_functions_0|redist5|delay_signals[0][20]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][20]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][20] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][20] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][21] (
	.clk(clk),
	.d(\fp_functions_0|redist5|delay_signals[0][21]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][21]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][21] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][21] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][22] (
	.clk(clk),
	.d(\fp_functions_0|redist5|delay_signals[0][22]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][22]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][22] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][22] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][23] (
	.clk(clk),
	.d(\fp_functions_0|redist5|delay_signals[0][23]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][23]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][23] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][23] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][24] (
	.clk(clk),
	.d(\fp_functions_0|redist5|delay_signals[0][24]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][24]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][24] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][24] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][25] (
	.clk(clk),
	.d(\fp_functions_0|redist5|delay_signals[0][25]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][25]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][25] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][25] .power_up = "low";

dffeas \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][26] (
	.clk(clk),
	.d(\fp_functions_0|redist5|delay_signals[0][26]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][26]~q ),
	.prn(vcc));
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][26] .is_wysiwyg = "true";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][26] .power_up = "low";

dffeas \fp_functions_0|redist15_inputreg|delay_signals[0][11] (
	.clk(clk),
	.d(\fp_functions_0|expSum_uid44_fpMulTest_o[11]~q ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist15_inputreg|delay_signals[0][11]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist15_inputreg|delay_signals[0][11] .is_wysiwyg = "true";
defparam \fp_functions_0|redist15_inputreg|delay_signals[0][11] .power_up = "low";

dffeas \fp_functions_0|redist6|delay_signals[0][0] (
	.clk(clk),
	.d(b[26]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist6|delay_signals[0][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist6|delay_signals[0][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist6|delay_signals[0][0] .power_up = "low";

dffeas \fp_functions_0|redist6|delay_signals[0][1] (
	.clk(clk),
	.d(b[27]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist6|delay_signals[0][1]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist6|delay_signals[0][1] .is_wysiwyg = "true";
defparam \fp_functions_0|redist6|delay_signals[0][1] .power_up = "low";

dffeas \fp_functions_0|redist6|delay_signals[0][2] (
	.clk(clk),
	.d(b[28]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist6|delay_signals[0][2]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist6|delay_signals[0][2] .is_wysiwyg = "true";
defparam \fp_functions_0|redist6|delay_signals[0][2] .power_up = "low";

dffeas \fp_functions_0|redist6|delay_signals[0][3] (
	.clk(clk),
	.d(b[29]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist6|delay_signals[0][3]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist6|delay_signals[0][3] .is_wysiwyg = "true";
defparam \fp_functions_0|redist6|delay_signals[0][3] .power_up = "low";

dffeas \fp_functions_0|redist6|delay_signals[0][4] (
	.clk(clk),
	.d(b[30]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist6|delay_signals[0][4]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist6|delay_signals[0][4] .is_wysiwyg = "true";
defparam \fp_functions_0|redist6|delay_signals[0][4] .power_up = "low";

dffeas \fp_functions_0|redist6|delay_signals[0][5] (
	.clk(clk),
	.d(b[31]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist6|delay_signals[0][5]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist6|delay_signals[0][5] .is_wysiwyg = "true";
defparam \fp_functions_0|redist6|delay_signals[0][5] .power_up = "low";

dffeas \fp_functions_0|redist6|delay_signals[0][6] (
	.clk(clk),
	.d(b[32]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist6|delay_signals[0][6]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist6|delay_signals[0][6] .is_wysiwyg = "true";
defparam \fp_functions_0|redist6|delay_signals[0][6] .power_up = "low";

dffeas \fp_functions_0|redist6|delay_signals[0][7] (
	.clk(clk),
	.d(b[33]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist6|delay_signals[0][7]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist6|delay_signals[0][7] .is_wysiwyg = "true";
defparam \fp_functions_0|redist6|delay_signals[0][7] .power_up = "low";

dffeas \fp_functions_0|redist6|delay_signals[0][8] (
	.clk(clk),
	.d(b[34]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist6|delay_signals[0][8]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist6|delay_signals[0][8] .is_wysiwyg = "true";
defparam \fp_functions_0|redist6|delay_signals[0][8] .power_up = "low";

dffeas \fp_functions_0|redist6|delay_signals[0][9] (
	.clk(clk),
	.d(b[35]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist6|delay_signals[0][9]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist6|delay_signals[0][9] .is_wysiwyg = "true";
defparam \fp_functions_0|redist6|delay_signals[0][9] .power_up = "low";

dffeas \fp_functions_0|redist6|delay_signals[0][10] (
	.clk(clk),
	.d(b[36]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist6|delay_signals[0][10]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist6|delay_signals[0][10] .is_wysiwyg = "true";
defparam \fp_functions_0|redist6|delay_signals[0][10] .power_up = "low";

dffeas \fp_functions_0|redist6|delay_signals[0][11] (
	.clk(clk),
	.d(b[37]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist6|delay_signals[0][11]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist6|delay_signals[0][11] .is_wysiwyg = "true";
defparam \fp_functions_0|redist6|delay_signals[0][11] .power_up = "low";

dffeas \fp_functions_0|redist6|delay_signals[0][12] (
	.clk(clk),
	.d(b[38]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist6|delay_signals[0][12]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist6|delay_signals[0][12] .is_wysiwyg = "true";
defparam \fp_functions_0|redist6|delay_signals[0][12] .power_up = "low";

dffeas \fp_functions_0|redist6|delay_signals[0][13] (
	.clk(clk),
	.d(b[39]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist6|delay_signals[0][13]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist6|delay_signals[0][13] .is_wysiwyg = "true";
defparam \fp_functions_0|redist6|delay_signals[0][13] .power_up = "low";

dffeas \fp_functions_0|redist6|delay_signals[0][14] (
	.clk(clk),
	.d(b[40]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist6|delay_signals[0][14]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist6|delay_signals[0][14] .is_wysiwyg = "true";
defparam \fp_functions_0|redist6|delay_signals[0][14] .power_up = "low";

dffeas \fp_functions_0|redist6|delay_signals[0][15] (
	.clk(clk),
	.d(b[41]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist6|delay_signals[0][15]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist6|delay_signals[0][15] .is_wysiwyg = "true";
defparam \fp_functions_0|redist6|delay_signals[0][15] .power_up = "low";

dffeas \fp_functions_0|redist6|delay_signals[0][16] (
	.clk(clk),
	.d(b[42]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist6|delay_signals[0][16]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist6|delay_signals[0][16] .is_wysiwyg = "true";
defparam \fp_functions_0|redist6|delay_signals[0][16] .power_up = "low";

dffeas \fp_functions_0|redist6|delay_signals[0][17] (
	.clk(clk),
	.d(b[43]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist6|delay_signals[0][17]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist6|delay_signals[0][17] .is_wysiwyg = "true";
defparam \fp_functions_0|redist6|delay_signals[0][17] .power_up = "low";

dffeas \fp_functions_0|redist6|delay_signals[0][18] (
	.clk(clk),
	.d(b[44]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist6|delay_signals[0][18]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist6|delay_signals[0][18] .is_wysiwyg = "true";
defparam \fp_functions_0|redist6|delay_signals[0][18] .power_up = "low";

dffeas \fp_functions_0|redist6|delay_signals[0][19] (
	.clk(clk),
	.d(b[45]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist6|delay_signals[0][19]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist6|delay_signals[0][19] .is_wysiwyg = "true";
defparam \fp_functions_0|redist6|delay_signals[0][19] .power_up = "low";

dffeas \fp_functions_0|redist6|delay_signals[0][20] (
	.clk(clk),
	.d(b[46]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist6|delay_signals[0][20]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist6|delay_signals[0][20] .is_wysiwyg = "true";
defparam \fp_functions_0|redist6|delay_signals[0][20] .power_up = "low";

dffeas \fp_functions_0|redist6|delay_signals[0][21] (
	.clk(clk),
	.d(b[47]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist6|delay_signals[0][21]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist6|delay_signals[0][21] .is_wysiwyg = "true";
defparam \fp_functions_0|redist6|delay_signals[0][21] .power_up = "low";

dffeas \fp_functions_0|redist6|delay_signals[0][22] (
	.clk(clk),
	.d(b[48]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist6|delay_signals[0][22]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist6|delay_signals[0][22] .is_wysiwyg = "true";
defparam \fp_functions_0|redist6|delay_signals[0][22] .power_up = "low";

dffeas \fp_functions_0|redist6|delay_signals[0][23] (
	.clk(clk),
	.d(b[49]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist6|delay_signals[0][23]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist6|delay_signals[0][23] .is_wysiwyg = "true";
defparam \fp_functions_0|redist6|delay_signals[0][23] .power_up = "low";

dffeas \fp_functions_0|redist6|delay_signals[0][24] (
	.clk(clk),
	.d(b[50]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist6|delay_signals[0][24]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist6|delay_signals[0][24] .is_wysiwyg = "true";
defparam \fp_functions_0|redist6|delay_signals[0][24] .power_up = "low";

dffeas \fp_functions_0|redist6|delay_signals[0][25] (
	.clk(clk),
	.d(b[51]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist6|delay_signals[0][25]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist6|delay_signals[0][25] .is_wysiwyg = "true";
defparam \fp_functions_0|redist6|delay_signals[0][25] .power_up = "low";

dffeas \fp_functions_0|redist6|delay_signals[0][26] (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist6|delay_signals[0][26]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist6|delay_signals[0][26] .is_wysiwyg = "true";
defparam \fp_functions_0|redist6|delay_signals[0][26] .power_up = "low";

dffeas \fp_functions_0|redist4|delay_signals[0][0] (
	.clk(clk),
	.d(a[0]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist4|delay_signals[0][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist4|delay_signals[0][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist4|delay_signals[0][0] .power_up = "low";

dffeas \fp_functions_0|redist4|delay_signals[0][1] (
	.clk(clk),
	.d(a[1]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist4|delay_signals[0][1]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist4|delay_signals[0][1] .is_wysiwyg = "true";
defparam \fp_functions_0|redist4|delay_signals[0][1] .power_up = "low";

dffeas \fp_functions_0|redist4|delay_signals[0][2] (
	.clk(clk),
	.d(a[2]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist4|delay_signals[0][2]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist4|delay_signals[0][2] .is_wysiwyg = "true";
defparam \fp_functions_0|redist4|delay_signals[0][2] .power_up = "low";

dffeas \fp_functions_0|redist4|delay_signals[0][3] (
	.clk(clk),
	.d(a[3]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist4|delay_signals[0][3]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist4|delay_signals[0][3] .is_wysiwyg = "true";
defparam \fp_functions_0|redist4|delay_signals[0][3] .power_up = "low";

dffeas \fp_functions_0|redist4|delay_signals[0][4] (
	.clk(clk),
	.d(a[4]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist4|delay_signals[0][4]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist4|delay_signals[0][4] .is_wysiwyg = "true";
defparam \fp_functions_0|redist4|delay_signals[0][4] .power_up = "low";

dffeas \fp_functions_0|redist4|delay_signals[0][5] (
	.clk(clk),
	.d(a[5]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist4|delay_signals[0][5]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist4|delay_signals[0][5] .is_wysiwyg = "true";
defparam \fp_functions_0|redist4|delay_signals[0][5] .power_up = "low";

dffeas \fp_functions_0|redist4|delay_signals[0][6] (
	.clk(clk),
	.d(a[6]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist4|delay_signals[0][6]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist4|delay_signals[0][6] .is_wysiwyg = "true";
defparam \fp_functions_0|redist4|delay_signals[0][6] .power_up = "low";

dffeas \fp_functions_0|redist4|delay_signals[0][7] (
	.clk(clk),
	.d(a[7]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist4|delay_signals[0][7]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist4|delay_signals[0][7] .is_wysiwyg = "true";
defparam \fp_functions_0|redist4|delay_signals[0][7] .power_up = "low";

dffeas \fp_functions_0|redist4|delay_signals[0][8] (
	.clk(clk),
	.d(a[8]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist4|delay_signals[0][8]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist4|delay_signals[0][8] .is_wysiwyg = "true";
defparam \fp_functions_0|redist4|delay_signals[0][8] .power_up = "low";

dffeas \fp_functions_0|redist4|delay_signals[0][9] (
	.clk(clk),
	.d(a[9]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist4|delay_signals[0][9]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist4|delay_signals[0][9] .is_wysiwyg = "true";
defparam \fp_functions_0|redist4|delay_signals[0][9] .power_up = "low";

dffeas \fp_functions_0|redist4|delay_signals[0][10] (
	.clk(clk),
	.d(a[10]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist4|delay_signals[0][10]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist4|delay_signals[0][10] .is_wysiwyg = "true";
defparam \fp_functions_0|redist4|delay_signals[0][10] .power_up = "low";

dffeas \fp_functions_0|redist4|delay_signals[0][11] (
	.clk(clk),
	.d(a[11]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist4|delay_signals[0][11]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist4|delay_signals[0][11] .is_wysiwyg = "true";
defparam \fp_functions_0|redist4|delay_signals[0][11] .power_up = "low";

dffeas \fp_functions_0|redist4|delay_signals[0][12] (
	.clk(clk),
	.d(a[12]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist4|delay_signals[0][12]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist4|delay_signals[0][12] .is_wysiwyg = "true";
defparam \fp_functions_0|redist4|delay_signals[0][12] .power_up = "low";

dffeas \fp_functions_0|redist4|delay_signals[0][13] (
	.clk(clk),
	.d(a[13]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist4|delay_signals[0][13]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist4|delay_signals[0][13] .is_wysiwyg = "true";
defparam \fp_functions_0|redist4|delay_signals[0][13] .power_up = "low";

dffeas \fp_functions_0|redist4|delay_signals[0][14] (
	.clk(clk),
	.d(a[14]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist4|delay_signals[0][14]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist4|delay_signals[0][14] .is_wysiwyg = "true";
defparam \fp_functions_0|redist4|delay_signals[0][14] .power_up = "low";

dffeas \fp_functions_0|redist4|delay_signals[0][15] (
	.clk(clk),
	.d(a[15]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist4|delay_signals[0][15]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist4|delay_signals[0][15] .is_wysiwyg = "true";
defparam \fp_functions_0|redist4|delay_signals[0][15] .power_up = "low";

dffeas \fp_functions_0|redist4|delay_signals[0][16] (
	.clk(clk),
	.d(a[16]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist4|delay_signals[0][16]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist4|delay_signals[0][16] .is_wysiwyg = "true";
defparam \fp_functions_0|redist4|delay_signals[0][16] .power_up = "low";

dffeas \fp_functions_0|redist4|delay_signals[0][17] (
	.clk(clk),
	.d(a[17]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist4|delay_signals[0][17]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist4|delay_signals[0][17] .is_wysiwyg = "true";
defparam \fp_functions_0|redist4|delay_signals[0][17] .power_up = "low";

dffeas \fp_functions_0|redist4|delay_signals[0][18] (
	.clk(clk),
	.d(a[18]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist4|delay_signals[0][18]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist4|delay_signals[0][18] .is_wysiwyg = "true";
defparam \fp_functions_0|redist4|delay_signals[0][18] .power_up = "low";

dffeas \fp_functions_0|redist4|delay_signals[0][19] (
	.clk(clk),
	.d(a[19]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist4|delay_signals[0][19]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist4|delay_signals[0][19] .is_wysiwyg = "true";
defparam \fp_functions_0|redist4|delay_signals[0][19] .power_up = "low";

dffeas \fp_functions_0|redist4|delay_signals[0][20] (
	.clk(clk),
	.d(a[20]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist4|delay_signals[0][20]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist4|delay_signals[0][20] .is_wysiwyg = "true";
defparam \fp_functions_0|redist4|delay_signals[0][20] .power_up = "low";

dffeas \fp_functions_0|redist4|delay_signals[0][21] (
	.clk(clk),
	.d(a[21]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist4|delay_signals[0][21]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist4|delay_signals[0][21] .is_wysiwyg = "true";
defparam \fp_functions_0|redist4|delay_signals[0][21] .power_up = "low";

dffeas \fp_functions_0|redist4|delay_signals[0][22] (
	.clk(clk),
	.d(a[22]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist4|delay_signals[0][22]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist4|delay_signals[0][22] .is_wysiwyg = "true";
defparam \fp_functions_0|redist4|delay_signals[0][22] .power_up = "low";

dffeas \fp_functions_0|redist4|delay_signals[0][23] (
	.clk(clk),
	.d(a[23]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist4|delay_signals[0][23]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist4|delay_signals[0][23] .is_wysiwyg = "true";
defparam \fp_functions_0|redist4|delay_signals[0][23] .power_up = "low";

dffeas \fp_functions_0|redist4|delay_signals[0][24] (
	.clk(clk),
	.d(a[24]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist4|delay_signals[0][24]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist4|delay_signals[0][24] .is_wysiwyg = "true";
defparam \fp_functions_0|redist4|delay_signals[0][24] .power_up = "low";

dffeas \fp_functions_0|redist4|delay_signals[0][25] (
	.clk(clk),
	.d(a[25]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist4|delay_signals[0][25]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist4|delay_signals[0][25] .is_wysiwyg = "true";
defparam \fp_functions_0|redist4|delay_signals[0][25] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][0] (
	.clk(clk),
	.d(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][0]~0_combout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][0] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][0] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][1] (
	.clk(clk),
	.d(b[0]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][1]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][1] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][1] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][2] (
	.clk(clk),
	.d(b[1]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][2]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][2] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][2] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][3] (
	.clk(clk),
	.d(b[2]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][3]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][3] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][3] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][4] (
	.clk(clk),
	.d(b[3]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][4]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][4] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][4] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][5] (
	.clk(clk),
	.d(b[4]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][5]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][5] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][5] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][6] (
	.clk(clk),
	.d(b[5]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][6]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][6] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][6] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][7] (
	.clk(clk),
	.d(b[6]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][7]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][7] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][7] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][8] (
	.clk(clk),
	.d(b[7]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][8]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][8] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][8] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][9] (
	.clk(clk),
	.d(b[8]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][9]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][9] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][9] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][10] (
	.clk(clk),
	.d(b[9]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][10]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][10] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][10] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][11] (
	.clk(clk),
	.d(b[10]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][11]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][11] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][11] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][12] (
	.clk(clk),
	.d(b[11]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][12]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][12] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][12] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][13] (
	.clk(clk),
	.d(b[12]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][13]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][13] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][13] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][14] (
	.clk(clk),
	.d(b[13]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][14]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][14] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][14] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][15] (
	.clk(clk),
	.d(b[14]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][15]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][15] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][15] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][16] (
	.clk(clk),
	.d(b[15]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][16]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][16] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][16] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][17] (
	.clk(clk),
	.d(b[16]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][17]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][17] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][17] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][18] (
	.clk(clk),
	.d(b[17]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][18]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][18] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][18] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][19] (
	.clk(clk),
	.d(b[18]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][19]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][19] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][19] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][20] (
	.clk(clk),
	.d(b[19]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][20]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][20] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][20] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][21] (
	.clk(clk),
	.d(b[20]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][21]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][21] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][21] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][22] (
	.clk(clk),
	.d(b[21]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][22]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][22] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][22] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][23] (
	.clk(clk),
	.d(b[22]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][23]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][23] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][23] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][24] (
	.clk(clk),
	.d(b[23]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][24]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][24] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][24] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][25] (
	.clk(clk),
	.d(b[24]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][25]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][25] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][25] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][26] (
	.clk(clk),
	.d(b[25]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][26]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][26] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][26] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][0] (
	.clk(clk),
	.d(a[26]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][0] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][0] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][1] (
	.clk(clk),
	.d(a[27]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][1]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][1] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][1] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][2] (
	.clk(clk),
	.d(a[28]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][2]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][2] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][2] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][3] (
	.clk(clk),
	.d(a[29]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][3]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][3] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][3] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][4] (
	.clk(clk),
	.d(a[30]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][4]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][4] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][4] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][5] (
	.clk(clk),
	.d(a[31]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][5]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][5] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][5] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][6] (
	.clk(clk),
	.d(a[32]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][6]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][6] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][6] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][7] (
	.clk(clk),
	.d(a[33]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][7]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][7] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][7] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][8] (
	.clk(clk),
	.d(a[34]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][8]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][8] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][8] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][9] (
	.clk(clk),
	.d(a[35]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][9]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][9] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][9] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][10] (
	.clk(clk),
	.d(a[36]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][10]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][10] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][10] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][11] (
	.clk(clk),
	.d(a[37]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][11]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][11] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][11] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][12] (
	.clk(clk),
	.d(a[38]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][12]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][12] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][12] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][13] (
	.clk(clk),
	.d(a[39]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][13]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][13] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][13] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][14] (
	.clk(clk),
	.d(a[40]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][14]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][14] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][14] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][15] (
	.clk(clk),
	.d(a[41]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][15]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][15] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][15] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][16] (
	.clk(clk),
	.d(a[42]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][16]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][16] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][16] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][17] (
	.clk(clk),
	.d(a[43]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][17]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][17] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][17] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][18] (
	.clk(clk),
	.d(a[44]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][18]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][18] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][18] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][19] (
	.clk(clk),
	.d(a[45]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][19]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][19] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][19] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][20] (
	.clk(clk),
	.d(a[46]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][20]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][20] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][20] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][21] (
	.clk(clk),
	.d(a[47]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][21]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][21] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][21] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][22] (
	.clk(clk),
	.d(a[48]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][22]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][22] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][22] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][23] (
	.clk(clk),
	.d(a[49]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][23]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][23] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][23] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][24] (
	.clk(clk),
	.d(a[50]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][24]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][24] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][24] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][25] (
	.clk(clk),
	.d(a[51]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][25]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][25] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][25] .power_up = "low";

dffeas \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][26] (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][26]~q ),
	.prn(vcc));
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][26] .is_wysiwyg = "true";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[1][26] .power_up = "low";

dffeas \fp_functions_0|redist7|delay_signals[0][0] (
	.clk(clk),
	.d(a[26]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist7|delay_signals[0][0]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist7|delay_signals[0][0] .is_wysiwyg = "true";
defparam \fp_functions_0|redist7|delay_signals[0][0] .power_up = "low";

dffeas \fp_functions_0|redist7|delay_signals[0][1] (
	.clk(clk),
	.d(a[27]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist7|delay_signals[0][1]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist7|delay_signals[0][1] .is_wysiwyg = "true";
defparam \fp_functions_0|redist7|delay_signals[0][1] .power_up = "low";

dffeas \fp_functions_0|redist7|delay_signals[0][2] (
	.clk(clk),
	.d(a[28]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist7|delay_signals[0][2]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist7|delay_signals[0][2] .is_wysiwyg = "true";
defparam \fp_functions_0|redist7|delay_signals[0][2] .power_up = "low";

dffeas \fp_functions_0|redist7|delay_signals[0][3] (
	.clk(clk),
	.d(a[29]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist7|delay_signals[0][3]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist7|delay_signals[0][3] .is_wysiwyg = "true";
defparam \fp_functions_0|redist7|delay_signals[0][3] .power_up = "low";

dffeas \fp_functions_0|redist7|delay_signals[0][4] (
	.clk(clk),
	.d(a[30]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist7|delay_signals[0][4]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist7|delay_signals[0][4] .is_wysiwyg = "true";
defparam \fp_functions_0|redist7|delay_signals[0][4] .power_up = "low";

dffeas \fp_functions_0|redist7|delay_signals[0][5] (
	.clk(clk),
	.d(a[31]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist7|delay_signals[0][5]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist7|delay_signals[0][5] .is_wysiwyg = "true";
defparam \fp_functions_0|redist7|delay_signals[0][5] .power_up = "low";

dffeas \fp_functions_0|redist7|delay_signals[0][6] (
	.clk(clk),
	.d(a[32]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist7|delay_signals[0][6]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist7|delay_signals[0][6] .is_wysiwyg = "true";
defparam \fp_functions_0|redist7|delay_signals[0][6] .power_up = "low";

dffeas \fp_functions_0|redist7|delay_signals[0][7] (
	.clk(clk),
	.d(a[33]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist7|delay_signals[0][7]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist7|delay_signals[0][7] .is_wysiwyg = "true";
defparam \fp_functions_0|redist7|delay_signals[0][7] .power_up = "low";

dffeas \fp_functions_0|redist7|delay_signals[0][8] (
	.clk(clk),
	.d(a[34]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist7|delay_signals[0][8]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist7|delay_signals[0][8] .is_wysiwyg = "true";
defparam \fp_functions_0|redist7|delay_signals[0][8] .power_up = "low";

dffeas \fp_functions_0|redist7|delay_signals[0][9] (
	.clk(clk),
	.d(a[35]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist7|delay_signals[0][9]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist7|delay_signals[0][9] .is_wysiwyg = "true";
defparam \fp_functions_0|redist7|delay_signals[0][9] .power_up = "low";

dffeas \fp_functions_0|redist7|delay_signals[0][10] (
	.clk(clk),
	.d(a[36]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist7|delay_signals[0][10]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist7|delay_signals[0][10] .is_wysiwyg = "true";
defparam \fp_functions_0|redist7|delay_signals[0][10] .power_up = "low";

dffeas \fp_functions_0|redist7|delay_signals[0][11] (
	.clk(clk),
	.d(a[37]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist7|delay_signals[0][11]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist7|delay_signals[0][11] .is_wysiwyg = "true";
defparam \fp_functions_0|redist7|delay_signals[0][11] .power_up = "low";

dffeas \fp_functions_0|redist7|delay_signals[0][12] (
	.clk(clk),
	.d(a[38]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist7|delay_signals[0][12]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist7|delay_signals[0][12] .is_wysiwyg = "true";
defparam \fp_functions_0|redist7|delay_signals[0][12] .power_up = "low";

dffeas \fp_functions_0|redist7|delay_signals[0][13] (
	.clk(clk),
	.d(a[39]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist7|delay_signals[0][13]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist7|delay_signals[0][13] .is_wysiwyg = "true";
defparam \fp_functions_0|redist7|delay_signals[0][13] .power_up = "low";

dffeas \fp_functions_0|redist7|delay_signals[0][14] (
	.clk(clk),
	.d(a[40]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist7|delay_signals[0][14]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist7|delay_signals[0][14] .is_wysiwyg = "true";
defparam \fp_functions_0|redist7|delay_signals[0][14] .power_up = "low";

dffeas \fp_functions_0|redist7|delay_signals[0][15] (
	.clk(clk),
	.d(a[41]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist7|delay_signals[0][15]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist7|delay_signals[0][15] .is_wysiwyg = "true";
defparam \fp_functions_0|redist7|delay_signals[0][15] .power_up = "low";

dffeas \fp_functions_0|redist7|delay_signals[0][16] (
	.clk(clk),
	.d(a[42]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist7|delay_signals[0][16]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist7|delay_signals[0][16] .is_wysiwyg = "true";
defparam \fp_functions_0|redist7|delay_signals[0][16] .power_up = "low";

dffeas \fp_functions_0|redist7|delay_signals[0][17] (
	.clk(clk),
	.d(a[43]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist7|delay_signals[0][17]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist7|delay_signals[0][17] .is_wysiwyg = "true";
defparam \fp_functions_0|redist7|delay_signals[0][17] .power_up = "low";

dffeas \fp_functions_0|redist7|delay_signals[0][18] (
	.clk(clk),
	.d(a[44]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist7|delay_signals[0][18]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist7|delay_signals[0][18] .is_wysiwyg = "true";
defparam \fp_functions_0|redist7|delay_signals[0][18] .power_up = "low";

dffeas \fp_functions_0|redist7|delay_signals[0][19] (
	.clk(clk),
	.d(a[45]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist7|delay_signals[0][19]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist7|delay_signals[0][19] .is_wysiwyg = "true";
defparam \fp_functions_0|redist7|delay_signals[0][19] .power_up = "low";

dffeas \fp_functions_0|redist7|delay_signals[0][20] (
	.clk(clk),
	.d(a[46]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist7|delay_signals[0][20]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist7|delay_signals[0][20] .is_wysiwyg = "true";
defparam \fp_functions_0|redist7|delay_signals[0][20] .power_up = "low";

dffeas \fp_functions_0|redist7|delay_signals[0][21] (
	.clk(clk),
	.d(a[47]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist7|delay_signals[0][21]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist7|delay_signals[0][21] .is_wysiwyg = "true";
defparam \fp_functions_0|redist7|delay_signals[0][21] .power_up = "low";

dffeas \fp_functions_0|redist7|delay_signals[0][22] (
	.clk(clk),
	.d(a[48]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist7|delay_signals[0][22]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist7|delay_signals[0][22] .is_wysiwyg = "true";
defparam \fp_functions_0|redist7|delay_signals[0][22] .power_up = "low";

dffeas \fp_functions_0|redist7|delay_signals[0][23] (
	.clk(clk),
	.d(a[49]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist7|delay_signals[0][23]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist7|delay_signals[0][23] .is_wysiwyg = "true";
defparam \fp_functions_0|redist7|delay_signals[0][23] .power_up = "low";

dffeas \fp_functions_0|redist7|delay_signals[0][24] (
	.clk(clk),
	.d(a[50]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist7|delay_signals[0][24]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist7|delay_signals[0][24] .is_wysiwyg = "true";
defparam \fp_functions_0|redist7|delay_signals[0][24] .power_up = "low";

dffeas \fp_functions_0|redist7|delay_signals[0][25] (
	.clk(clk),
	.d(a[51]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist7|delay_signals[0][25]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist7|delay_signals[0][25] .is_wysiwyg = "true";
defparam \fp_functions_0|redist7|delay_signals[0][25] .power_up = "low";

dffeas \fp_functions_0|redist7|delay_signals[0][26] (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist7|delay_signals[0][26]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist7|delay_signals[0][26] .is_wysiwyg = "true";
defparam \fp_functions_0|redist7|delay_signals[0][26] .power_up = "low";

dffeas \fp_functions_0|redist5|delay_signals[0][1] (
	.clk(clk),
	.d(b[0]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist5|delay_signals[0][1]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist5|delay_signals[0][1] .is_wysiwyg = "true";
defparam \fp_functions_0|redist5|delay_signals[0][1] .power_up = "low";

dffeas \fp_functions_0|redist5|delay_signals[0][2] (
	.clk(clk),
	.d(b[1]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist5|delay_signals[0][2]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist5|delay_signals[0][2] .is_wysiwyg = "true";
defparam \fp_functions_0|redist5|delay_signals[0][2] .power_up = "low";

dffeas \fp_functions_0|redist5|delay_signals[0][3] (
	.clk(clk),
	.d(b[2]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist5|delay_signals[0][3]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist5|delay_signals[0][3] .is_wysiwyg = "true";
defparam \fp_functions_0|redist5|delay_signals[0][3] .power_up = "low";

dffeas \fp_functions_0|redist5|delay_signals[0][4] (
	.clk(clk),
	.d(b[3]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist5|delay_signals[0][4]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist5|delay_signals[0][4] .is_wysiwyg = "true";
defparam \fp_functions_0|redist5|delay_signals[0][4] .power_up = "low";

dffeas \fp_functions_0|redist5|delay_signals[0][5] (
	.clk(clk),
	.d(b[4]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist5|delay_signals[0][5]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist5|delay_signals[0][5] .is_wysiwyg = "true";
defparam \fp_functions_0|redist5|delay_signals[0][5] .power_up = "low";

dffeas \fp_functions_0|redist5|delay_signals[0][6] (
	.clk(clk),
	.d(b[5]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist5|delay_signals[0][6]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist5|delay_signals[0][6] .is_wysiwyg = "true";
defparam \fp_functions_0|redist5|delay_signals[0][6] .power_up = "low";

dffeas \fp_functions_0|redist5|delay_signals[0][7] (
	.clk(clk),
	.d(b[6]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist5|delay_signals[0][7]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist5|delay_signals[0][7] .is_wysiwyg = "true";
defparam \fp_functions_0|redist5|delay_signals[0][7] .power_up = "low";

dffeas \fp_functions_0|redist5|delay_signals[0][8] (
	.clk(clk),
	.d(b[7]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist5|delay_signals[0][8]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist5|delay_signals[0][8] .is_wysiwyg = "true";
defparam \fp_functions_0|redist5|delay_signals[0][8] .power_up = "low";

dffeas \fp_functions_0|redist5|delay_signals[0][9] (
	.clk(clk),
	.d(b[8]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist5|delay_signals[0][9]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist5|delay_signals[0][9] .is_wysiwyg = "true";
defparam \fp_functions_0|redist5|delay_signals[0][9] .power_up = "low";

dffeas \fp_functions_0|redist5|delay_signals[0][10] (
	.clk(clk),
	.d(b[9]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist5|delay_signals[0][10]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist5|delay_signals[0][10] .is_wysiwyg = "true";
defparam \fp_functions_0|redist5|delay_signals[0][10] .power_up = "low";

dffeas \fp_functions_0|redist5|delay_signals[0][11] (
	.clk(clk),
	.d(b[10]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist5|delay_signals[0][11]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist5|delay_signals[0][11] .is_wysiwyg = "true";
defparam \fp_functions_0|redist5|delay_signals[0][11] .power_up = "low";

dffeas \fp_functions_0|redist5|delay_signals[0][12] (
	.clk(clk),
	.d(b[11]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist5|delay_signals[0][12]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist5|delay_signals[0][12] .is_wysiwyg = "true";
defparam \fp_functions_0|redist5|delay_signals[0][12] .power_up = "low";

dffeas \fp_functions_0|redist5|delay_signals[0][13] (
	.clk(clk),
	.d(b[12]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist5|delay_signals[0][13]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist5|delay_signals[0][13] .is_wysiwyg = "true";
defparam \fp_functions_0|redist5|delay_signals[0][13] .power_up = "low";

dffeas \fp_functions_0|redist5|delay_signals[0][14] (
	.clk(clk),
	.d(b[13]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist5|delay_signals[0][14]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist5|delay_signals[0][14] .is_wysiwyg = "true";
defparam \fp_functions_0|redist5|delay_signals[0][14] .power_up = "low";

dffeas \fp_functions_0|redist5|delay_signals[0][15] (
	.clk(clk),
	.d(b[14]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist5|delay_signals[0][15]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist5|delay_signals[0][15] .is_wysiwyg = "true";
defparam \fp_functions_0|redist5|delay_signals[0][15] .power_up = "low";

dffeas \fp_functions_0|redist5|delay_signals[0][16] (
	.clk(clk),
	.d(b[15]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist5|delay_signals[0][16]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist5|delay_signals[0][16] .is_wysiwyg = "true";
defparam \fp_functions_0|redist5|delay_signals[0][16] .power_up = "low";

dffeas \fp_functions_0|redist5|delay_signals[0][17] (
	.clk(clk),
	.d(b[16]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist5|delay_signals[0][17]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist5|delay_signals[0][17] .is_wysiwyg = "true";
defparam \fp_functions_0|redist5|delay_signals[0][17] .power_up = "low";

dffeas \fp_functions_0|redist5|delay_signals[0][18] (
	.clk(clk),
	.d(b[17]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist5|delay_signals[0][18]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist5|delay_signals[0][18] .is_wysiwyg = "true";
defparam \fp_functions_0|redist5|delay_signals[0][18] .power_up = "low";

dffeas \fp_functions_0|redist5|delay_signals[0][19] (
	.clk(clk),
	.d(b[18]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist5|delay_signals[0][19]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist5|delay_signals[0][19] .is_wysiwyg = "true";
defparam \fp_functions_0|redist5|delay_signals[0][19] .power_up = "low";

dffeas \fp_functions_0|redist5|delay_signals[0][20] (
	.clk(clk),
	.d(b[19]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist5|delay_signals[0][20]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist5|delay_signals[0][20] .is_wysiwyg = "true";
defparam \fp_functions_0|redist5|delay_signals[0][20] .power_up = "low";

dffeas \fp_functions_0|redist5|delay_signals[0][21] (
	.clk(clk),
	.d(b[20]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist5|delay_signals[0][21]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist5|delay_signals[0][21] .is_wysiwyg = "true";
defparam \fp_functions_0|redist5|delay_signals[0][21] .power_up = "low";

dffeas \fp_functions_0|redist5|delay_signals[0][22] (
	.clk(clk),
	.d(b[21]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist5|delay_signals[0][22]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist5|delay_signals[0][22] .is_wysiwyg = "true";
defparam \fp_functions_0|redist5|delay_signals[0][22] .power_up = "low";

dffeas \fp_functions_0|redist5|delay_signals[0][23] (
	.clk(clk),
	.d(b[22]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist5|delay_signals[0][23]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist5|delay_signals[0][23] .is_wysiwyg = "true";
defparam \fp_functions_0|redist5|delay_signals[0][23] .power_up = "low";

dffeas \fp_functions_0|redist5|delay_signals[0][24] (
	.clk(clk),
	.d(b[23]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist5|delay_signals[0][24]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist5|delay_signals[0][24] .is_wysiwyg = "true";
defparam \fp_functions_0|redist5|delay_signals[0][24] .power_up = "low";

dffeas \fp_functions_0|redist5|delay_signals[0][25] (
	.clk(clk),
	.d(b[24]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist5|delay_signals[0][25]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist5|delay_signals[0][25] .is_wysiwyg = "true";
defparam \fp_functions_0|redist5|delay_signals[0][25] .power_up = "low";

dffeas \fp_functions_0|redist5|delay_signals[0][26] (
	.clk(clk),
	.d(b[25]),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|redist5|delay_signals[0][26]~q ),
	.prn(vcc));
defparam \fp_functions_0|redist5|delay_signals[0][26] .is_wysiwyg = "true";
defparam \fp_functions_0|redist5|delay_signals[0][26] .power_up = "low";

dffeas \fp_functions_0|expSum_uid44_fpMulTest_o[11] (
	.clk(clk),
	.d(\fp_functions_0|add_4~45_sumout ),
	.asdata(vcc),
	.clrn(!areset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(en[0]),
	.q(\fp_functions_0|expSum_uid44_fpMulTest_o[11]~q ),
	.prn(vcc));
defparam \fp_functions_0|expSum_uid44_fpMulTest_o[11] .is_wysiwyg = "true";
defparam \fp_functions_0|expSum_uid44_fpMulTest_o[11] .power_up = "low";

twentynm_lcell_comb \fp_functions_0|reduce_nor_7~11 (
	.dataa(!\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[1]~q ),
	.datab(!\fp_functions_0|fracRPostNorm_uid53_fpMulTest_q[0]~q ),
	.datac(!\fp_functions_0|redist12|delay_signals[0][29]~q ),
	.datad(!\fp_functions_0|redist12|delay_signals[0][35]~q ),
	.datae(!\fp_functions_0|redist12|delay_signals[0][17]~q ),
	.dataf(!\fp_functions_0|redist12|delay_signals[0][23]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|reduce_nor_7~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|reduce_nor_7~11 .extended_lut = "off";
defparam \fp_functions_0|reduce_nor_7~11 .lut_mask = 64'h2000000000000000;
defparam \fp_functions_0|reduce_nor_7~11 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|reduce_nor_7~12 (
	.dataa(!\fp_functions_0|reduce_nor_7~5_combout ),
	.datab(!\fp_functions_0|reduce_nor_7~6_combout ),
	.datac(!\fp_functions_0|reduce_nor_7~7_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|reduce_nor_7~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|reduce_nor_7~12 .extended_lut = "off";
defparam \fp_functions_0|reduce_nor_7~12 .lut_mask = 64'h0101010101010101;
defparam \fp_functions_0|reduce_nor_7~12 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|redist11|delay_signals[0][53]~0 (
	.dataa(!\fp_functions_0|redist15_outputreg|delay_signals[0][0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|redist11|delay_signals[0][53]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|redist11|delay_signals[0][53]~0 .extended_lut = "off";
defparam \fp_functions_0|redist11|delay_signals[0][53]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \fp_functions_0|redist11|delay_signals[0][53]~0 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][0]~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][0]~0 .extended_lut = "off";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][0]~0 .lut_mask = 64'h0000000000000000;
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_c0[0][0]~0 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][0]~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][0]~0 .extended_lut = "off";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][0]~0 .lut_mask = 64'h0000000000000000;
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_a0[0][0]~0 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][0]~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][0]~0 .extended_lut = "off";
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][0]~0 .lut_mask = 64'h0000000000000000;
defparam \fp_functions_0|sm0_uid128_prod_uid47_fpMulTest_cma_c0[0][0]~0 .shared_arith = "off";

twentynm_lcell_comb \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][0]~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][0]~0 .extended_lut = "off";
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][0]~0 .lut_mask = 64'h0000000000000000;
defparam \fp_functions_0|multSumOfTwoTS_uid118_prod_uid47_fpMulTest_cma_a0[1][0]~0 .shared_arith = "off";

assign q[0] = \fp_functions_0|Mux_64~0_combout ;

assign q[1] = \fp_functions_0|Mux_63~0_combout ;

assign q[2] = \fp_functions_0|Mux_62~0_combout ;

assign q[3] = \fp_functions_0|Mux_61~0_combout ;

assign q[4] = \fp_functions_0|Mux_60~0_combout ;

assign q[5] = \fp_functions_0|Mux_59~0_combout ;

assign q[6] = \fp_functions_0|Mux_58~0_combout ;

assign q[7] = \fp_functions_0|Mux_57~0_combout ;

assign q[8] = \fp_functions_0|Mux_56~0_combout ;

assign q[9] = \fp_functions_0|Mux_55~0_combout ;

assign q[10] = \fp_functions_0|Mux_54~0_combout ;

assign q[11] = \fp_functions_0|Mux_53~0_combout ;

assign q[12] = \fp_functions_0|Mux_52~0_combout ;

assign q[13] = \fp_functions_0|Mux_51~0_combout ;

assign q[14] = \fp_functions_0|Mux_50~0_combout ;

assign q[15] = \fp_functions_0|Mux_49~0_combout ;

assign q[16] = \fp_functions_0|Mux_48~0_combout ;

assign q[17] = \fp_functions_0|Mux_47~0_combout ;

assign q[18] = \fp_functions_0|Mux_46~0_combout ;

assign q[19] = \fp_functions_0|Mux_45~0_combout ;

assign q[20] = \fp_functions_0|Mux_44~0_combout ;

assign q[21] = \fp_functions_0|Mux_43~0_combout ;

assign q[22] = \fp_functions_0|Mux_42~0_combout ;

assign q[23] = \fp_functions_0|Mux_41~0_combout ;

assign q[24] = \fp_functions_0|Mux_40~0_combout ;

assign q[25] = \fp_functions_0|Mux_39~0_combout ;

assign q[26] = \fp_functions_0|Mux_38~0_combout ;

assign q[27] = \fp_functions_0|Mux_37~0_combout ;

assign q[28] = \fp_functions_0|Mux_36~0_combout ;

assign q[29] = \fp_functions_0|Mux_35~0_combout ;

assign q[30] = \fp_functions_0|Mux_34~0_combout ;

assign q[31] = \fp_functions_0|Mux_33~0_combout ;

assign q[32] = \fp_functions_0|Mux_32~0_combout ;

assign q[33] = \fp_functions_0|Mux_31~0_combout ;

assign q[34] = \fp_functions_0|Mux_30~0_combout ;

assign q[35] = \fp_functions_0|Mux_29~0_combout ;

assign q[36] = \fp_functions_0|Mux_28~0_combout ;

assign q[37] = \fp_functions_0|Mux_27~0_combout ;

assign q[38] = \fp_functions_0|Mux_26~0_combout ;

assign q[39] = \fp_functions_0|Mux_25~0_combout ;

assign q[40] = \fp_functions_0|Mux_24~0_combout ;

assign q[41] = \fp_functions_0|Mux_23~0_combout ;

assign q[42] = \fp_functions_0|Mux_22~0_combout ;

assign q[43] = \fp_functions_0|Mux_21~0_combout ;

assign q[44] = \fp_functions_0|Mux_20~0_combout ;

assign q[45] = \fp_functions_0|Mux_19~0_combout ;

assign q[46] = \fp_functions_0|Mux_18~0_combout ;

assign q[47] = \fp_functions_0|Mux_17~0_combout ;

assign q[48] = \fp_functions_0|Mux_16~0_combout ;

assign q[49] = \fp_functions_0|Mux_15~0_combout ;

assign q[50] = \fp_functions_0|Mux_14~0_combout ;

assign q[51] = \fp_functions_0|Mux_13~0_combout ;

assign q[52] = \fp_functions_0|Mux_12~0_combout ;

assign q[53] = \fp_functions_0|Mux_12~1_combout ;

assign q[54] = \fp_functions_0|Mux_12~2_combout ;

assign q[55] = \fp_functions_0|Mux_12~3_combout ;

assign q[56] = \fp_functions_0|Mux_12~4_combout ;

assign q[57] = \fp_functions_0|Mux_12~5_combout ;

assign q[58] = \fp_functions_0|Mux_12~6_combout ;

assign q[59] = \fp_functions_0|Mux_12~7_combout ;

assign q[60] = \fp_functions_0|Mux_12~8_combout ;

assign q[61] = \fp_functions_0|Mux_12~9_combout ;

assign q[62] = \fp_functions_0|Mux_12~10_combout ;

assign q[63] = \fp_functions_0|i1071~combout ;

endmodule
