-- ram32x64.vhd

-- Generated using ACDS version 16.0 211

library IEEE;
--library ram_1port_160;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity ram32x64 is
	port (
		data    : in  std_logic_vector(63 downto 0) := (others => '0'); --  ram_input.datain
		address : in  std_logic_vector(4 downto 0)  := (others => '0'); --           .address
		wren    : in  std_logic                     := '0';             --           .wren
		clock   : in  std_logic                     := '0';             --           .clk
		q       : out std_logic_vector(63 downto 0)                     -- ram_output.dataout
	);
end entity ram32x64;

architecture rtl of ram32x64 is
	component ram32x64_ram_1port_160_lcifr2i is
		port (
			data    : in  std_logic_vector(63 downto 0) := (others => 'X'); -- datain
			address : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- address
			wren    : in  std_logic                     := 'X';             -- wren
			clock   : in  std_logic                     := 'X';             -- clk
			q       : out std_logic_vector(63 downto 0)                     -- dataout
		);
	end component ram32x64_ram_1port_160_lcifr2i;

--	for ram_1port_0 : ram32x64_ram_1port_160_lcifr2i
--		use entity ram_1port_160.ram32x64_ram_1port_160_lcifr2i;
begin

	ram_1port_0 : component ram32x64_ram_1port_160_lcifr2i
		port map (
			data    => data,    --  ram_input.datain
			address => address, --           .address
			wren    => wren,    --           .wren
			clock   => clock,   --           .clk
			q       => q        -- ram_output.dataout
		);

end architecture rtl; -- of ram32x64
